module ASCIIRenderer (
  input [10:0] x, y,
  input [7:0] ascii,
  output reg hit
);

reg [10:0] pixel_x, pixel_y;

always @ (ascii or x or y)
begin
  pixel_x = (ascii - 33) + x;
  pixel_y = y;
end

always @ (*)
if((pixel_x >= 52 && pixel_x < 54 && pixel_y >= 1 && pixel_y < 24) || (pixel_x >= 19 && pixel_x < 21 && pixel_y >= 2 && pixel_y < 9) || (pixel_x >= 24 && pixel_x < 26 && pixel_y >= 2 && pixel_y < 9) || (pixel_x >= 73 && pixel_x < 75 && pixel_y == 2) || (pixel_x == 81 && pixel_y >= 2 && pixel_y < 4) || (pixel_x >= 96 && pixel_x < 99 && pixel_y >= 2 && pixel_y < 9) || (pixel_x >= 115 && pixel_x < 118 && pixel_y >= 2 && pixel_y < 4) || (pixel_x >= 122 && pixel_x < 125 && pixel_y >= 2 && pixel_y < 4) || (pixel_x == 142 && pixel_y >= 2 && pixel_y < 14) || (pixel_x == 223 && pixel_y >= 2 && pixel_y < 4) || (pixel_x == 232 && pixel_y >= 2 && pixel_y < 4) || (pixel_x == 262 && pixel_y >= 2 && pixel_y < 4) || (pixel_x == 276 && pixel_y >= 2 && pixel_y < 4) || (pixel_x >= 323 && pixel_x < 325 && pixel_y >= 2 && pixel_y < 4) || (pixel_x == 352 && pixel_y >= 2 && pixel_y < 4) || (pixel_x == 367 && pixel_y >= 2 && pixel_y < 5) || (pixel_x >= 456 && pixel_x < 458 && pixel_y >= 2 && pixel_y < 4) || (pixel_x == 472 && pixel_y >= 2 && pixel_y < 4) || (pixel_x == 519 && pixel_y >= 2 && pixel_y < 4) || (pixel_x == 579 && pixel_y >= 2 && pixel_y < 4) || (pixel_x == 697 && pixel_y >= 2 && pixel_y < 4) || (pixel_x == 727 && pixel_y >= 2 && pixel_y < 4) || (pixel_x >= 757 && pixel_x < 759 && pixel_y >= 2 && pixel_y < 4) || (pixel_x >= 874 && pixel_x < 877 && pixel_y >= 2 && pixel_y < 26) || (pixel_x >= 877 && pixel_x < 884 && pixel_y >= 2 && pixel_y < 4) || (pixel_x >= 886 && pixel_x < 888 && pixel_y >= 2 && pixel_y < 4) || (pixel_x >= 901 && pixel_x < 911 && pixel_y >= 2 && pixel_y < 4) || (pixel_x >= 950 && pixel_x < 952 && pixel_y >= 2 && pixel_y < 4) || (pixel_x >= 977 && pixel_x < 979 && pixel_y >= 2 && pixel_y < 22) || (pixel_x >= 1016 && pixel_x < 1018 && pixel_y >= 2 && pixel_y < 22) || (pixel_x >= 1043 && pixel_x < 1049 && pixel_y >= 2 && pixel_y < 4) || (pixel_x >= 1067 && pixel_x < 1069 && pixel_y >= 2 && pixel_y < 22) || (pixel_x >= 1086 && pixel_x < 1088 && pixel_y >= 2 && pixel_y < 5) || (pixel_x >= 1104 && pixel_x < 1106 && pixel_y >= 2 && pixel_y < 5) || (pixel_x >= 1113 && pixel_x < 1115 && pixel_y >= 2 && pixel_y < 22) || (pixel_x >= 1127 && pixel_x < 1133 && pixel_y >= 2 && pixel_y < 4) || (pixel_x >= 1358 && pixel_x < 1364 && pixel_y >= 2 && pixel_y < 4) || (pixel_x == 1372 && pixel_y >= 2 && pixel_y < 23) || (pixel_x >= 1382 && pixel_x < 1387 && pixel_y >= 2 && pixel_y < 4) || (pixel_x >= 6 && pixel_x < 9 && pixel_y >= 3 && pixel_y < 13) || (pixel_x == 18 && pixel_y == 3) || (pixel_x == 26 && pixel_y == 3) || (pixel_x >= 36 && pixel_x < 38 && pixel_y >= 3 && pixel_y < 6) || (pixel_x == 42 && pixel_y >= 3 && pixel_y < 7) || (pixel_x >= 50 && pixel_x < 52 && pixel_y >= 3 && pixel_y < 5) || (pixel_x >= 54 && pixel_x < 57 && pixel_y >= 3 && pixel_y < 5) || (pixel_x >= 62 && pixel_x < 66 && pixel_y >= 3 && pixel_y < 5) || (pixel_x >= 72 && pixel_x < 74 && pixel_y >= 3 && pixel_y < 5) || (pixel_x >= 78 && pixel_x < 80 && pixel_y >= 3 && pixel_y < 5) || (pixel_x == 80 && pixel_y == 3) || (pixel_x >= 82 && pixel_x < 84 && pixel_y >= 3 && pixel_y < 5) || (pixel_x >= 113 && pixel_x < 115 && pixel_y >= 3 && pixel_y < 5) || (pixel_x >= 125 && pixel_x < 127 && pixel_y >= 3 && pixel_y < 5) || (pixel_x == 141 && pixel_y >= 3 && pixel_y < 14) || (pixel_x == 143 && pixel_y >= 3 && pixel_y < 14) || (pixel_x == 222 && pixel_y >= 3 && pixel_y < 6) || (pixel_x >= 229 && pixel_x < 232 && pixel_y >= 3 && pixel_y < 5) || (pixel_x >= 233 && pixel_x < 236 && pixel_y >= 3 && pixel_y < 5) || (pixel_x >= 246 && pixel_x < 249 && pixel_y >= 3 && pixel_y < 6) || (pixel_x >= 258 && pixel_x < 261 && pixel_y >= 3 && pixel_y < 5) || (pixel_x == 261 && pixel_y == 3) || (pixel_x >= 263 && pixel_x < 266 && pixel_y >= 3 && pixel_y < 5) || (pixel_x >= 272 && pixel_x < 275 && pixel_y >= 3 && pixel_y < 5) || (pixel_x == 275 && pixel_y == 3) || (pixel_x >= 277 && pixel_x < 281 && pixel_y == 3) || (pixel_x >= 293 && pixel_x < 296 && pixel_y >= 3 && pixel_y < 8) || (pixel_x >= 302 && pixel_x < 305 && pixel_y >= 3 && pixel_y < 12) || (pixel_x >= 305 && pixel_x < 313 && pixel_y >= 3 && pixel_y < 5) || (pixel_x >= 320 && pixel_x < 323 && pixel_y >= 3 && pixel_y < 5) || (pixel_x >= 325 && pixel_x < 328 && pixel_y >= 3 && pixel_y < 5) || (pixel_x >= 332 && pixel_x < 344 && pixel_y >= 3 && pixel_y < 5) || (pixel_x >= 350 && pixel_x < 352 && pixel_y >= 3 && pixel_y < 5) || (pixel_x >= 353 && pixel_x < 356 && pixel_y >= 3 && pixel_y < 5) || (pixel_x >= 364 && pixel_x < 367 && pixel_y >= 3 && pixel_y < 5) || (pixel_x >= 368 && pixel_x < 371 && pixel_y >= 3 && pixel_y < 5) || (pixel_x >= 453 && pixel_x < 456 && pixel_y >= 3 && pixel_y < 5) || (pixel_x >= 458 && pixel_x < 461 && pixel_y == 3) || (pixel_x >= 469 && pixel_x < 472 && pixel_y == 3) || (pixel_x >= 473 && pixel_x < 477 && pixel_y == 3) || (pixel_x >= 486 && pixel_x < 489 && pixel_y >= 3 && pixel_y < 8) || (pixel_x >= 497 && pixel_x < 500 && pixel_y >= 3 && pixel_y < 22) || (pixel_x >= 500 && pixel_x < 505 && pixel_y >= 3 && pixel_y < 5) || (pixel_x >= 516 && pixel_x < 519 && pixel_y >= 3 && pixel_y < 5) || (pixel_x >= 520 && pixel_x < 523 && pixel_y == 3) || (pixel_x >= 527 && pixel_x < 535 && pixel_y >= 3 && pixel_y < 5) || (pixel_x >= 543 && pixel_x < 553 && pixel_y >= 3 && pixel_y < 5) || (pixel_x >= 558 && pixel_x < 568 && pixel_y >= 3 && pixel_y < 5) || (pixel_x >= 576 && pixel_x < 579 && pixel_y >= 3 && pixel_y < 5) || (pixel_x >= 580 && pixel_x < 583 && pixel_y == 3) || (pixel_x >= 587 && pixel_x < 589 && pixel_y >= 3 && pixel_y < 22) || (pixel_x >= 596 && pixel_x < 599 && pixel_y >= 3 && pixel_y < 22) || (pixel_x >= 602 && pixel_x < 613 && pixel_y >= 3 && pixel_y < 5) || (pixel_x >= 620 && pixel_x < 627 && pixel_y >= 3 && pixel_y < 5) || (pixel_x >= 632 && pixel_x < 634 && pixel_y >= 3 && pixel_y < 22) || (pixel_x >= 641 && pixel_x < 643 && pixel_y >= 3 && pixel_y < 5) || (pixel_x == 643 && pixel_y == 3) || (pixel_x >= 648 && pixel_x < 650 && pixel_y >= 3 && pixel_y < 22) || (pixel_x >= 661 && pixel_x < 663 && pixel_y >= 3 && pixel_y < 22) || (pixel_x >= 672 && pixel_x < 674 && pixel_y >= 3 && pixel_y < 22) || (pixel_x >= 677 && pixel_x < 679 && pixel_y >= 3 && pixel_y < 22) || (pixel_x >= 686 && pixel_x < 689 && pixel_y >= 3 && pixel_y < 22) || (pixel_x >= 694 && pixel_x < 697 && pixel_y >= 3 && pixel_y < 5) || (pixel_x >= 698 && pixel_x < 701 && pixel_y == 3) || (pixel_x >= 707 && pixel_x < 710 && pixel_y >= 3 && pixel_y < 22) || (pixel_x >= 710 && pixel_x < 716 && pixel_y >= 3 && pixel_y < 5) || (pixel_x >= 724 && pixel_x < 727 && pixel_y >= 3 && pixel_y < 5) || (pixel_x >= 728 && pixel_x < 731 && pixel_y == 3) || (pixel_x >= 737 && pixel_x < 746 && pixel_y >= 3 && pixel_y < 5) || (pixel_x >= 754 && pixel_x < 757 && pixel_y >= 3 && pixel_y < 5) || (pixel_x >= 759 && pixel_x < 762 && pixel_y == 3) || (pixel_x >= 766 && pixel_x < 780 && pixel_y >= 3 && pixel_y < 5) || (pixel_x >= 782 && pixel_x < 784 && pixel_y >= 3 && pixel_y < 20) || (pixel_x >= 791 && pixel_x < 794 && pixel_y >= 3 && pixel_y < 17) || (pixel_x >= 796 && pixel_x < 798 && pixel_y >= 3 && pixel_y < 6) || (pixel_x >= 807 && pixel_x < 809 && pixel_y >= 3 && pixel_y < 7) || (pixel_x == 809 && pixel_y == 3) || (pixel_x >= 811 && pixel_x < 813 && pixel_y >= 3 && pixel_y < 12) || (pixel_x >= 816 && pixel_x < 819 && pixel_y >= 3 && pixel_y < 9) || (pixel_x >= 823 && pixel_x < 825 && pixel_y >= 3 && pixel_y < 5) || (pixel_x >= 827 && pixel_x < 829 && pixel_y >= 3 && pixel_y < 5) || (pixel_x >= 836 && pixel_x < 838 && pixel_y >= 3 && pixel_y < 6) || (pixel_x == 838 && pixel_y == 3) || (pixel_x >= 841 && pixel_x < 844 && pixel_y == 3) || (pixel_x >= 852 && pixel_x < 854 && pixel_y >= 3 && pixel_y < 5) || (pixel_x >= 857 && pixel_x < 868 && pixel_y >= 3 && pixel_y < 5) || (pixel_x == 922 && pixel_y >= 3 && pixel_y < 8) || (pixel_x == 952 && pixel_y >= 3 && pixel_y < 6) || (pixel_x == 1042 && pixel_y >= 3 && pixel_y < 22) || (pixel_x == 1106 && pixel_y == 3) || (pixel_x == 1357 && pixel_y >= 3 && pixel_y < 14) || (pixel_x == 1373 && pixel_y >= 3 && pixel_y < 22) || (pixel_x == 1387 && pixel_y >= 3 && pixel_y < 14) || (pixel_x == 41 && pixel_y >= 4 && pixel_y < 11) || (pixel_x == 49 && pixel_y >= 4 && pixel_y < 12) || (pixel_x == 61 && pixel_y >= 4 && pixel_y < 12) || (pixel_x == 66 && pixel_y >= 4 && pixel_y < 16) || (pixel_x == 77 && pixel_y >= 4 && pixel_y < 10) || (pixel_x == 84 && pixel_y >= 4 && pixel_y < 7) || (pixel_x == 112 && pixel_y >= 4 && pixel_y < 7) || (pixel_x == 127 && pixel_y >= 4 && pixel_y < 7) || (pixel_x == 221 && pixel_y >= 4 && pixel_y < 8) || (pixel_x == 228 && pixel_y >= 4 && pixel_y < 10) || (pixel_x == 236 && pixel_y >= 4 && pixel_y < 10) || (pixel_x == 245 && pixel_y >= 4 && pixel_y < 7) || (pixel_x == 257 && pixel_y >= 4 && pixel_y < 6) || (pixel_x == 266 && pixel_y >= 4 && pixel_y < 10) || (pixel_x >= 278 && pixel_x < 282 && pixel_y == 4) || (pixel_x == 319 && pixel_y >= 4 && pixel_y < 8) || (pixel_x == 349 && pixel_y >= 4 && pixel_y < 11) || (pixel_x == 356 && pixel_y >= 4 && pixel_y < 10) || (pixel_x == 363 && pixel_y >= 4 && pixel_y < 8) || (pixel_x == 371 && pixel_y >= 4 && pixel_y < 20) || (pixel_x >= 459 && pixel_x < 462 && pixel_y == 4) || (pixel_x >= 468 && pixel_x < 470 && pixel_y == 4) || (pixel_x >= 475 && pixel_x < 478 && pixel_y == 4) || (pixel_x == 505 && pixel_y >= 4 && pixel_y < 11) || (pixel_x >= 514 && pixel_x < 516 && pixel_y >= 4 && pixel_y < 7) || (pixel_x >= 521 && pixel_x < 523 && pixel_y == 4) || (pixel_x >= 535 && pixel_x < 537 && pixel_y >= 4 && pixel_y < 7) || (pixel_x >= 574 && pixel_x < 576 && pixel_y >= 4 && pixel_y < 7) || (pixel_x >= 581 && pixel_x < 583 && pixel_y == 4) || (pixel_x == 640 && pixel_y >= 4 && pixel_y < 8) || (pixel_x == 663 && pixel_y >= 4 && pixel_y < 11) || (pixel_x == 679 && pixel_y >= 4 && pixel_y < 9) || (pixel_x == 693 && pixel_y >= 4 && pixel_y < 11) || (pixel_x >= 699 && pixel_x < 702 && pixel_y == 4) || (pixel_x == 716 && pixel_y >= 4 && pixel_y < 14) || (pixel_x == 723 && pixel_y >= 4 && pixel_y < 11) || (pixel_x >= 729 && pixel_x < 732 && pixel_y == 4) || (pixel_x == 746 && pixel_y >= 4 && pixel_y < 11) || (pixel_x == 753 && pixel_y >= 4 && pixel_y < 11) || (pixel_x >= 760 && pixel_x < 762 && pixel_y == 4) || (pixel_x == 798 && pixel_y >= 4 && pixel_y < 13) || (pixel_x == 829 && pixel_y >= 4 && pixel_y < 9) || (pixel_x >= 842 && pixel_x < 844 && pixel_y >= 4 && pixel_y < 6) || (pixel_x == 851 && pixel_y >= 4 && pixel_y < 9) || (pixel_x >= 887 && pixel_x < 889 && pixel_y >= 4 && pixel_y < 6) || (pixel_x >= 909 && pixel_x < 911 && pixel_y >= 4 && pixel_y < 27) || (pixel_x == 951 && pixel_y == 4) || (pixel_x == 953 && pixel_y >= 4 && pixel_y < 6) || (pixel_x == 1041 && pixel_y >= 4 && pixel_y < 22) || (pixel_x == 1043 && pixel_y == 4) || (pixel_x >= 1131 && pixel_x < 1133 && pixel_y >= 4 && pixel_y < 22) || (pixel_x >= 1250 && pixel_x < 1252 && pixel_y >= 4 && pixel_y < 20) || (pixel_x == 1358 && pixel_y >= 4 && pixel_y < 13) || (pixel_x == 1386 && pixel_y == 4) || (pixel_x == 1388 && pixel_y >= 4 && pixel_y < 8) || (pixel_x == 48 && pixel_y >= 5 && pixel_y < 11) || (pixel_x == 50 && pixel_y == 5) || (pixel_x == 56 && pixel_y == 5) || (pixel_x == 60 && pixel_y >= 5 && pixel_y < 10) || (pixel_x == 62 && pixel_y == 5) || (pixel_x == 65 && pixel_y >= 5 && pixel_y < 7) || (pixel_x >= 71 && pixel_x < 73 && pixel_y == 5) || (pixel_x == 78 && pixel_y >= 5 && pixel_y < 14) || (pixel_x == 83 && pixel_y >= 5 && pixel_y < 9) || (pixel_x == 111 && pixel_y >= 5 && pixel_y < 8) || (pixel_x == 113 && pixel_y == 5) || (pixel_x == 126 && pixel_y == 5) || (pixel_x == 128 && pixel_y >= 5 && pixel_y < 8) || (pixel_x >= 137 && pixel_x < 140 && pixel_y >= 5 && pixel_y < 7) || (pixel_x >= 145 && pixel_x < 148 && pixel_y >= 5 && pixel_y < 7) || (pixel_x == 227 && pixel_y >= 5 && pixel_y < 20) || (pixel_x == 229 && pixel_y >= 5 && pixel_y < 7) || (pixel_x == 235 && pixel_y >= 5 && pixel_y < 10) || (pixel_x == 237 && pixel_y >= 5 && pixel_y < 20) || (pixel_x >= 243 && pixel_x < 245 && pixel_y >= 5 && pixel_y < 7) || (pixel_x == 265 && pixel_y >= 5 && pixel_y < 11) || (pixel_x == 267 && pixel_y >= 5 && pixel_y < 8) || (pixel_x >= 279 && pixel_x < 282 && pixel_y == 5) || (pixel_x == 292 && pixel_y >= 5 && pixel_y < 8) || (pixel_x == 318 && pixel_y >= 5 && pixel_y < 21) || (pixel_x == 320 && pixel_y == 5) || (pixel_x >= 341 && pixel_x < 344 && pixel_y >= 5 && pixel_y < 7) || (pixel_x == 348 && pixel_y >= 5 && pixel_y < 10) || (pixel_x == 350 && pixel_y == 5) || (pixel_x == 355 && pixel_y >= 5 && pixel_y < 11) || (pixel_x == 357 && pixel_y >= 5 && pixel_y < 8) || (pixel_x == 362 && pixel_y >= 5 && pixel_y < 13) || (pixel_x == 364 && pixel_y == 5) || (pixel_x >= 369 && pixel_x < 371 && pixel_y == 5) || (pixel_x >= 460 && pixel_x < 463 && pixel_y >= 5 && pixel_y < 8) || (pixel_x >= 467 && pixel_x < 469 && pixel_y == 5) || (pixel_x >= 477 && pixel_x < 479 && pixel_y >= 5 && pixel_y < 7) || (pixel_x == 489 && pixel_y >= 5 && pixel_y < 14) || (pixel_x == 504 && pixel_y == 5) || (pixel_x == 506 && pixel_y >= 5 && pixel_y < 11) || (pixel_x == 513 && pixel_y >= 5 && pixel_y < 20) || (pixel_x == 516 && pixel_y == 5) || (pixel_x >= 527 && pixel_x < 529 && pixel_y >= 5 && pixel_y < 22) || (pixel_x == 534 && pixel_y == 5) || (pixel_x >= 543 && pixel_x < 545 && pixel_y >= 5 && pixel_y < 22) || (pixel_x >= 558 && pixel_x < 560 && pixel_y >= 5 && pixel_y < 22) || (pixel_x == 573 && pixel_y >= 5 && pixel_y < 20) || (pixel_x == 576 && pixel_y == 5) || (pixel_x >= 606 && pixel_x < 609 && pixel_y >= 5 && pixel_y < 22) || (pixel_x >= 624 && pixel_x < 627 && pixel_y >= 5 && pixel_y < 19) || (pixel_x == 641 && pixel_y >= 5 && pixel_y < 7) || (pixel_x == 671 && pixel_y >= 5 && pixel_y < 10) || (pixel_x == 692 && pixel_y >= 5 && pixel_y < 20) || (pixel_x == 694 && pixel_y >= 5 && pixel_y < 7) || (pixel_x >= 700 && pixel_x < 703 && pixel_y == 5) || (pixel_x == 715 && pixel_y == 5) || (pixel_x == 717 && pixel_y >= 5 && pixel_y < 13) || (pixel_x == 722 && pixel_y >= 5 && pixel_y < 19) || (pixel_x == 724 && pixel_y >= 5 && pixel_y < 7) || (pixel_x >= 730 && pixel_x < 733 && pixel_y == 5) || (pixel_x >= 737 && pixel_x < 739 && pixel_y >= 5 && pixel_y < 22) || (pixel_x >= 744 && pixel_x < 746 && pixel_y == 5) || (pixel_x == 747 && pixel_y >= 5 && pixel_y < 10) || (pixel_x >= 754 && pixel_x < 756 && pixel_y == 5) || (pixel_x >= 771 && pixel_x < 774 && pixel_y >= 5 && pixel_y < 22) || (pixel_x == 823 && pixel_y >= 5 && pixel_y < 14) || (pixel_x == 828 && pixel_y >= 5 && pixel_y < 7) || (pixel_x == 835 && pixel_y >= 5 && pixel_y < 9) || (pixel_x == 844 && pixel_y >= 5 && pixel_y < 10) || (pixel_x == 852 && pixel_y >= 5 && pixel_y < 7) || (pixel_x >= 865 && pixel_x < 868 && pixel_y >= 5 && pixel_y < 7) || (pixel_x == 889 && pixel_y >= 5 && pixel_y < 9) || (pixel_x == 921 && pixel_y >= 5 && pixel_y < 9) || (pixel_x == 923 && pixel_y >= 5 && pixel_y < 9) || (pixel_x == 954 && pixel_y == 5) || (pixel_x == 36 && pixel_y >= 6 && pixel_y < 10) || (pixel_x == 47 && pixel_y >= 6 && pixel_y < 10) || (pixel_x == 67 && pixel_y >= 6 && pixel_y < 9) || (pixel_x >= 70 && pixel_x < 72 && pixel_y >= 6 && pixel_y < 8) || (pixel_x == 76 && pixel_y == 6) || (pixel_x == 110 && pixel_y >= 6 && pixel_y < 10) || (pixel_x == 129 && pixel_y >= 6 && pixel_y < 10) || (pixel_x == 140 && pixel_y >= 6 && pixel_y < 10) || (pixel_x == 144 && pixel_y >= 6 && pixel_y < 10) || (pixel_x == 220 && pixel_y >= 6 && pixel_y < 9) || (pixel_x == 242 && pixel_y >= 6 && pixel_y < 8) || (pixel_x >= 247 && pixel_x < 249 && pixel_y >= 6 && pixel_y < 22) || (pixel_x >= 280 && pixel_x < 282 && pixel_y >= 6 && pixel_y < 10) || (pixel_x == 291 && pixel_y >= 6 && pixel_y < 10) || (pixel_x == 361 && pixel_y >= 6 && pixel_y < 12) || (pixel_x == 370 && pixel_y >= 6 && pixel_y < 8) || (pixel_x == 372 && pixel_y >= 6 && pixel_y < 19) || (pixel_x >= 466 && pixel_x < 468 && pixel_y >= 6 && pixel_y < 8) || (pixel_x == 485 && pixel_y >= 6 && pixel_y < 13) || (pixel_x == 537 && pixel_y >= 6 && pixel_y < 19) || (pixel_x == 639 && pixel_y >= 6 && pixel_y < 9) || (pixel_x == 680 && pixel_y >= 6 && pixel_y < 11) || (pixel_x >= 701 && pixel_x < 703 && pixel_y >= 6 && pixel_y < 9) || (pixel_x == 718 && pixel_y >= 6 && pixel_y < 11) || (pixel_x >= 731 && pixel_x < 733 && pixel_y >= 6 && pixel_y < 9) || (pixel_x == 745 && pixel_y == 6) || (pixel_x == 752 && pixel_y >= 6 && pixel_y < 9) || (pixel_x == 754 && pixel_y >= 6 && pixel_y < 12) || (pixel_x == 797 && pixel_y >= 6 && pixel_y < 9) || (pixel_x == 806 && pixel_y >= 6 && pixel_y < 14) || (pixel_x == 822 && pixel_y >= 6 && pixel_y < 22) || (pixel_x == 830 && pixel_y >= 6 && pixel_y < 11) || (pixel_x == 834 && pixel_y >= 6 && pixel_y < 11) || (pixel_x == 836 && pixel_y == 6) || (pixel_x == 843 && pixel_y >= 6 && pixel_y < 8) || (pixel_x == 845 && pixel_y >= 6 && pixel_y < 12) || (pixel_x == 850 && pixel_y >= 6 && pixel_y < 10) || (pixel_x == 888 && pixel_y >= 6 && pixel_y < 8) || (pixel_x == 1040 && pixel_y >= 6 && pixel_y < 22) || (pixel_x == 1386 && pixel_y >= 6 && pixel_y < 13) || (pixel_x == 35 && pixel_y >= 7 && pixel_y < 13) || (pixel_x == 82 && pixel_y >= 7 && pixel_y < 10) || (pixel_x == 109 && pixel_y >= 7 && pixel_y < 22) || (pixel_x == 130 && pixel_y >= 7 && pixel_y < 22) || (pixel_x == 139 && pixel_y == 7) || (pixel_x == 145 && pixel_y == 7) || (pixel_x == 219 && pixel_y >= 7 && pixel_y < 11) || (pixel_x == 238 && pixel_y >= 7 && pixel_y < 18) || (pixel_x == 243 && pixel_y == 7) || (pixel_x == 317 && pixel_y >= 7 && pixel_y < 19) || (pixel_x >= 341 && pixel_x < 343 && pixel_y == 7) || (pixel_x >= 471 && pixel_x < 476 && pixel_y >= 7 && pixel_y < 9) || (pixel_x == 478 && pixel_y >= 7 && pixel_y < 10) || (pixel_x == 507 && pixel_y == 7) || (pixel_x == 512 && pixel_y >= 7 && pixel_y < 18) || (pixel_x == 514 && pixel_y >= 7 && pixel_y < 9) || (pixel_x == 536 && pixel_y >= 7 && pixel_y < 10) || (pixel_x == 572 && pixel_y >= 7 && pixel_y < 18) || (pixel_x == 574 && pixel_y >= 7 && pixel_y < 9) || (pixel_x == 638 && pixel_y >= 7 && pixel_y < 11) || (pixel_x == 664 && pixel_y >= 7 && pixel_y < 13) || (pixel_x == 670 && pixel_y >= 7 && pixel_y < 13) || (pixel_x == 703 && pixel_y >= 7 && pixel_y < 18) || (pixel_x == 733 && pixel_y >= 7 && pixel_y < 18) || (pixel_x == 799 && pixel_y >= 7 && pixel_y < 16) || (pixel_x == 807 && pixel_y >= 7 && pixel_y < 10) || (pixel_x == 819 && pixel_y >= 7 && pixel_y < 18) || (pixel_x == 831 && pixel_y >= 7 && pixel_y < 16) || (pixel_x == 849 && pixel_y >= 7 && pixel_y < 12) || (pixel_x >= 864 && pixel_x < 866 && pixel_y >= 7 && pixel_y < 10) || (pixel_x == 866 && pixel_y == 7) || (pixel_x == 890 && pixel_y >= 7 && pixel_y < 11) || (pixel_x == 920 && pixel_y >= 7 && pixel_y < 12) || (pixel_x == 924 && pixel_y >= 7 && pixel_y < 11) || (pixel_x >= 31 && pixel_x < 35 && pixel_y >= 8 && pixel_y < 10) || (pixel_x >= 37 && pixel_x < 41 && pixel_y >= 8 && pixel_y < 10) || (pixel_x >= 42 && pixel_x < 44 && pixel_y >= 8 && pixel_y < 10) || (pixel_x >= 69 && pixel_x < 71 && pixel_y >= 8 && pixel_y < 10) || (pixel_x == 226 && pixel_y >= 8 && pixel_y < 17) || (pixel_x == 234 && pixel_y >= 8 && pixel_y < 11) || (pixel_x == 279 && pixel_y >= 8 && pixel_y < 14) || (pixel_x == 290 && pixel_y >= 8 && pixel_y < 11) || (pixel_x >= 294 && pixel_x < 296 && pixel_y >= 8 && pixel_y < 22) || (pixel_x >= 340 && pixel_x < 342 && pixel_y >= 8 && pixel_y < 10) || (pixel_x == 350 && pixel_y >= 8 && pixel_y < 15) || (pixel_x >= 381 && pixel_x < 384 && pixel_y >= 8 && pixel_y < 11) || (pixel_x >= 396 && pixel_x < 399 && pixel_y >= 8 && pixel_y < 11) || (pixel_x >= 459 && pixel_x < 462 && pixel_y >= 8 && pixel_y < 10) || (pixel_x == 466 && pixel_y >= 8 && pixel_y < 19) || (pixel_x >= 469 && pixel_x < 471 && pixel_y >= 8 && pixel_y < 10) || (pixel_x == 479 && pixel_y >= 8 && pixel_y < 14) || (pixel_x == 486 && pixel_y >= 8 && pixel_y < 10) || (pixel_x == 488 && pixel_y >= 8 && pixel_y < 10) || (pixel_x == 490 && pixel_y >= 8 && pixel_y < 18) || (pixel_x == 538 && pixel_y >= 8 && pixel_y < 17) || (pixel_x == 637 && pixel_y >= 8 && pixel_y < 16) || (pixel_x == 681 && pixel_y >= 8 && pixel_y < 13) || (pixel_x == 691 && pixel_y >= 8 && pixel_y < 17) || (pixel_x == 721 && pixel_y >= 8 && pixel_y < 17) || (pixel_x == 833 && pixel_y >= 8 && pixel_y < 16) || (pixel_x == 846 && pixel_y >= 8 && pixel_y < 22) || (pixel_x == 863 && pixel_y >= 8 && pixel_y < 13) || (pixel_x >= 966 && pixel_x < 973 && pixel_y >= 8 && pixel_y < 10) || (pixel_x >= 983 && pixel_x < 986 && pixel_y >= 8 && pixel_y < 10) || (pixel_x >= 996 && pixel_x < 1003 && pixel_y >= 8 && pixel_y < 10) || (pixel_x >= 1011 && pixel_x < 1016 && pixel_y >= 8 && pixel_y < 10) || (pixel_x >= 1026 && pixel_x < 1031 && pixel_y >= 8 && pixel_y < 10) || (pixel_x >= 1056 && pixel_x < 1063 && pixel_y >= 8 && pixel_y < 10) || (pixel_x >= 1073 && pixel_x < 1076 && pixel_y >= 8 && pixel_y < 10) || (pixel_x >= 1082 && pixel_x < 1088 && pixel_y >= 8 && pixel_y < 10) || (pixel_x >= 1099 && pixel_x < 1106 && pixel_y >= 8 && pixel_y < 10) || (pixel_x >= 1121 && pixel_x < 1123 && pixel_y >= 8 && pixel_y < 10) || (pixel_x == 1123 && pixel_y == 8) || (pixel_x >= 1141 && pixel_x < 1143 && pixel_y >= 8 && pixel_y < 22) || (pixel_x >= 1145 && pixel_x < 1148 && pixel_y >= 8 && pixel_y < 11) || (pixel_x >= 1151 && pixel_x < 1153 && pixel_y >= 8 && pixel_y < 10) || (pixel_x >= 1157 && pixel_x < 1159 && pixel_y >= 8 && pixel_y < 22) || (pixel_x >= 1163 && pixel_x < 1166 && pixel_y >= 8 && pixel_y < 10) || (pixel_x >= 1175 && pixel_x < 1180 && pixel_y >= 8 && pixel_y < 10) || (pixel_x >= 1187 && pixel_x < 1189 && pixel_y >= 8 && pixel_y < 27) || (pixel_x >= 1193 && pixel_x < 1196 && pixel_y >= 8 && pixel_y < 10) || (pixel_x >= 1206 && pixel_x < 1213 && pixel_y >= 8 && pixel_y < 10) || (pixel_x >= 1218 && pixel_x < 1220 && pixel_y >= 8 && pixel_y < 22) || (pixel_x >= 1224 && pixel_x < 1228 && pixel_y >= 8 && pixel_y < 10) || (pixel_x >= 1235 && pixel_x < 1242 && pixel_y >= 8 && pixel_y < 10) || (pixel_x >= 1262 && pixel_x < 1264 && pixel_y >= 8 && pixel_y < 20) || (pixel_x >= 1271 && pixel_x < 1273 && pixel_y >= 8 && pixel_y < 22) || (pixel_x >= 1276 && pixel_x < 1278 && pixel_y >= 8 && pixel_y < 10) || (pixel_x >= 1288 && pixel_x < 1290 && pixel_y == 8) || (pixel_x == 1291 && pixel_y >= 8 && pixel_y < 15) || (pixel_x >= 1297 && pixel_x < 1299 && pixel_y >= 8 && pixel_y < 13) || (pixel_x >= 1303 && pixel_x < 1305 && pixel_y >= 8 && pixel_y < 11) || (pixel_x >= 1307 && pixel_x < 1309 && pixel_y >= 8 && pixel_y < 10) || (pixel_x >= 1316 && pixel_x < 1318 && pixel_y >= 8 && pixel_y < 10) || (pixel_x >= 1321 && pixel_x < 1323 && pixel_y >= 8 && pixel_y < 10) || (pixel_x >= 1333 && pixel_x < 1335 && pixel_y == 8) || (pixel_x >= 1337 && pixel_x < 1348 && pixel_y >= 8 && pixel_y < 10) || (pixel_x == 50 && pixel_y >= 9 && pixel_y < 12) || (pixel_x == 65 && pixel_y >= 9 && pixel_y < 12) || (pixel_x == 68 && pixel_y >= 9 && pixel_y < 21) || (pixel_x >= 79 && pixel_x < 82 && pixel_y >= 9 && pixel_y < 13) || (pixel_x == 97 && pixel_y == 9) || (pixel_x == 108 && pixel_y >= 9 && pixel_y < 20) || (pixel_x == 131 && pixel_y >= 9 && pixel_y < 20) || (pixel_x >= 138 && pixel_x < 140 && pixel_y >= 9 && pixel_y < 11) || (pixel_x >= 145 && pixel_x < 147 && pixel_y >= 9 && pixel_y < 11) || (pixel_x == 157 && pixel_y >= 9 && pixel_y < 22) || (pixel_x == 218 && pixel_y >= 9 && pixel_y < 13) || (pixel_x == 233 && pixel_y >= 9 && pixel_y < 13) || (pixel_x == 264 && pixel_y >= 9 && pixel_y < 13) || (pixel_x == 289 && pixel_y >= 9 && pixel_y < 13) || (pixel_x == 339 && pixel_y >= 9 && pixel_y < 12) || (pixel_x == 351 && pixel_y >= 9 && pixel_y < 14) || (pixel_x == 354 && pixel_y >= 9 && pixel_y < 15) || (pixel_x == 373 && pixel_y >= 9 && pixel_y < 16) || (pixel_x == 418 && pixel_y >= 9 && pixel_y < 11) || (pixel_x >= 436 && pixel_x < 438 && pixel_y >= 9 && pixel_y < 11) || (pixel_x == 465 && pixel_y >= 9 && pixel_y < 16) || (pixel_x >= 474 && pixel_x < 476 && pixel_y >= 9 && pixel_y < 16) || (pixel_x == 484 && pixel_y >= 9 && pixel_y < 18) || (pixel_x == 665 && pixel_y >= 9 && pixel_y < 16) || (pixel_x == 702 && pixel_y >= 9 && pixel_y < 20) || (pixel_x == 732 && pixel_y >= 9 && pixel_y < 20) || (pixel_x == 745 && pixel_y >= 9 && pixel_y < 12) || (pixel_x == 755 && pixel_y >= 9 && pixel_y < 12) || (pixel_x == 805 && pixel_y >= 9 && pixel_y < 17) || (pixel_x >= 815 && pixel_x < 817 && pixel_y >= 9 && pixel_y < 13) || (pixel_x == 818 && pixel_y >= 9 && pixel_y < 13) || (pixel_x == 832 && pixel_y >= 9 && pixel_y < 15) || (pixel_x == 848 && pixel_y >= 9 && pixel_y < 22) || (pixel_x == 891 && pixel_y >= 9 && pixel_y < 13) || (pixel_x == 919 && pixel_y >= 9 && pixel_y < 14) || (pixel_x == 925 && pixel_y >= 9 && pixel_y < 13) || (pixel_x >= 964 && pixel_x < 966 && pixel_y >= 9 && pixel_y < 11) || (pixel_x >= 981 && pixel_x < 983 && pixel_y >= 9 && pixel_y < 11) || (pixel_x == 986 && pixel_y >= 9 && pixel_y < 20) || (pixel_x == 995 && pixel_y >= 9 && pixel_y < 12) || (pixel_x == 1003 && pixel_y >= 9 && pixel_y < 11) || (pixel_x >= 1009 && pixel_x < 1011 && pixel_y >= 9 && pixel_y < 12) || (pixel_x >= 1024 && pixel_x < 1026 && pixel_y >= 9 && pixel_y < 11) || (pixel_x == 1031 && pixel_y >= 9 && pixel_y < 16) || (pixel_x >= 1037 && pixel_x < 1040 && pixel_y >= 9 && pixel_y < 11) || (pixel_x >= 1043 && pixel_x < 1048 && pixel_y >= 9 && pixel_y < 11) || (pixel_x >= 1054 && pixel_x < 1056 && pixel_y >= 9 && pixel_y < 12) || (pixel_x >= 1071 && pixel_x < 1073 && pixel_y >= 9 && pixel_y < 11) || (pixel_x == 1076 && pixel_y >= 9 && pixel_y < 22) || (pixel_x == 1098 && pixel_y == 9) || (pixel_x == 1120 && pixel_y >= 9 && pixel_y < 12) || (pixel_x == 1144 && pixel_y >= 9 && pixel_y < 11) || (pixel_x == 1150 && pixel_y >= 9 && pixel_y < 11) || (pixel_x == 1153 && pixel_y >= 9 && pixel_y < 22) || (pixel_x >= 1161 && pixel_x < 1163 && pixel_y >= 9 && pixel_y < 11) || (pixel_x == 1166 && pixel_y >= 9 && pixel_y < 22) || (pixel_x >= 1173 && pixel_x < 1175 && pixel_y >= 9 && pixel_y < 12) || (pixel_x >= 1180 && pixel_x < 1182 && pixel_y >= 9 && pixel_y < 11) || (pixel_x >= 1191 && pixel_x < 1193 && pixel_y >= 9 && pixel_y < 11) || (pixel_x >= 1196 && pixel_x < 1198 && pixel_y >= 9 && pixel_y < 19) || (pixel_x == 1205 && pixel_y >= 9 && pixel_y < 12) || (pixel_x == 1220 && pixel_y >= 9 && pixel_y < 22) || (pixel_x >= 1222 && pixel_x < 1224 && pixel_y >= 9 && pixel_y < 11) || (pixel_x >= 1233 && pixel_x < 1235 && pixel_y >= 9 && pixel_y < 14) || (pixel_x >= 1247 && pixel_x < 1250 && pixel_y >= 9 && pixel_y < 11) || (pixel_x >= 1252 && pixel_x < 1258 && pixel_y >= 9 && pixel_y < 11) || (pixel_x == 1278 && pixel_y >= 9 && pixel_y < 15) || (pixel_x >= 1287 && pixel_x < 1289 && pixel_y >= 9 && pixel_y < 11) || (pixel_x == 1292 && pixel_y >= 9 && pixel_y < 21) || (pixel_x == 1296 && pixel_y >= 9 && pixel_y < 16) || (pixel_x == 1309 && pixel_y >= 9 && pixel_y < 13) || (pixel_x == 1315 && pixel_y >= 9 && pixel_y < 13) || (pixel_x == 1323 && pixel_y >= 9 && pixel_y < 14) || (pixel_x >= 1332 && pixel_x < 1334 && pixel_y >= 9 && pixel_y < 12) || (pixel_x == 34 && pixel_y >= 10 && pixel_y < 17) || (pixel_x == 40 && pixel_y >= 10 && pixel_y < 14) || (pixel_x == 51 && pixel_y >= 10 && pixel_y < 13) || (pixel_x == 62 && pixel_y >= 10 && pixel_y < 12) || (pixel_x == 64 && pixel_y >= 10 && pixel_y < 12) || (pixel_x == 67 && pixel_y >= 10 && pixel_y < 15) || (pixel_x == 69 && pixel_y == 10) || (pixel_x == 137 && pixel_y == 10) || (pixel_x == 147 && pixel_y == 10) || (pixel_x >= 277 && pixel_x < 279 && pixel_y >= 10 && pixel_y < 13) || (pixel_x == 280 && pixel_y == 10) || (pixel_x == 288 && pixel_y >= 10 && pixel_y < 14) || (pixel_x >= 305 && pixel_x < 309 && pixel_y >= 10 && pixel_y < 12) || (pixel_x == 316 && pixel_y >= 10 && pixel_y < 16) || (pixel_x >= 322 && pixel_x < 325 && pixel_y >= 10 && pixel_y < 12) || (pixel_x == 338 && pixel_y >= 10 && pixel_y < 14) || (pixel_x == 340 && pixel_y == 10) || (pixel_x >= 352 && pixel_x < 354 && pixel_y >= 10 && pixel_y < 13) || (pixel_x == 370 && pixel_y >= 10 && pixel_y < 13) || (pixel_x >= 416 && pixel_x < 418 && pixel_y >= 10 && pixel_y < 12) || (pixel_x >= 438 && pixel_x < 440 && pixel_y >= 10 && pixel_y < 12) || (pixel_x >= 458 && pixel_x < 460 && pixel_y >= 10 && pixel_y < 12) || (pixel_x == 460 && pixel_y == 10) || (pixel_x >= 468 && pixel_x < 470 && pixel_y >= 10 && pixel_y < 15) || (pixel_x == 504 && pixel_y >= 10 && pixel_y < 15) || (pixel_x == 636 && pixel_y >= 10 && pixel_y < 15) || (pixel_x == 669 && pixel_y >= 10 && pixel_y < 16) || (pixel_x == 682 && pixel_y >= 10 && pixel_y < 15) || (pixel_x == 756 && pixel_y >= 10 && pixel_y < 13) || (pixel_x == 813 && pixel_y >= 10 && pixel_y < 22) || (pixel_x == 847 && pixel_y >= 10 && pixel_y < 22) || (pixel_x == 862 && pixel_y >= 10 && pixel_y < 15) || (pixel_x == 864 && pixel_y >= 10 && pixel_y < 12) || (pixel_x == 892 && pixel_y >= 10 && pixel_y < 14) || (pixel_x == 963 && pixel_y >= 10 && pixel_y < 22) || (pixel_x == 966 && pixel_y == 10) || (pixel_x >= 971 && pixel_x < 973 && pixel_y >= 10 && pixel_y < 22) || (pixel_x >= 979 && pixel_x < 981 && pixel_y >= 10 && pixel_y < 12) || (pixel_x >= 984 && pixel_x < 986 && pixel_y == 10) || (pixel_x == 987 && pixel_y >= 10 && pixel_y < 19) || (pixel_x == 994 && pixel_y >= 10 && pixel_y < 21) || (pixel_x == 996 && pixel_y == 10) || (pixel_x == 1002 && pixel_y == 10) || (pixel_x == 1008 && pixel_y >= 10 && pixel_y < 21) || (pixel_x == 1011 && pixel_y == 10) || (pixel_x == 1023 && pixel_y >= 10 && pixel_y < 20) || (pixel_x == 1026 && pixel_y == 10) || (pixel_x == 1030 && pixel_y == 10) || (pixel_x == 1032 && pixel_y >= 10 && pixel_y < 16) || (pixel_x == 1053 && pixel_y >= 10 && pixel_y < 21) || (pixel_x == 1056 && pixel_y == 10) || (pixel_x >= 1061 && pixel_x < 1063 && pixel_y >= 10 && pixel_y < 25) || (pixel_x >= 1069 && pixel_x < 1071 && pixel_y >= 10 && pixel_y < 12) || (pixel_x == 1075 && pixel_y == 10) || (pixel_x == 1077 && pixel_y >= 10 && pixel_y < 22) || (pixel_x >= 1086 && pixel_x < 1088 && pixel_y >= 10 && pixel_y < 22) || (pixel_x >= 1104 && pixel_x < 1106 && pixel_y >= 10 && pixel_y < 25) || (pixel_x == 1119 && pixel_y >= 10 && pixel_y < 13) || (pixel_x == 1121 && pixel_y == 10) || (pixel_x == 1143 && pixel_y >= 10 && pixel_y < 13) || (pixel_x >= 1148 && pixel_x < 1150 && pixel_y >= 10 && pixel_y < 12) || (pixel_x == 1152 && pixel_y >= 10 && pixel_y < 22) || (pixel_x >= 1159 && pixel_x < 1161 && pixel_y >= 10 && pixel_y < 12) || (pixel_x == 1165 && pixel_y == 10) || (pixel_x == 1167 && pixel_y >= 10 && pixel_y < 22) || (pixel_x == 1175 && pixel_y == 10) || (pixel_x == 1182 && pixel_y >= 10 && pixel_y < 20) || (pixel_x == 1190 && pixel_y >= 10 && pixel_y < 12) || (pixel_x >= 1194 && pixel_x < 1196 && pixel_y == 10) || (pixel_x == 1204 && pixel_y >= 10 && pixel_y < 13) || (pixel_x == 1206 && pixel_y == 10) || (pixel_x >= 1211 && pixel_x < 1213 && pixel_y >= 10 && pixel_y < 27) || (pixel_x == 1221 && pixel_y >= 10 && pixel_y < 13) || (pixel_x >= 1226 && pixel_x < 1228 && pixel_y >= 10 && pixel_y < 13) || (pixel_x == 1235 && pixel_y == 10) || (pixel_x == 1246 && pixel_y == 10) || (pixel_x == 1277 && pixel_y >= 10 && pixel_y < 13) || (pixel_x == 1308 && pixel_y == 10) || (pixel_x == 1310 && pixel_y >= 10 && pixel_y < 14) || (pixel_x == 1314 && pixel_y >= 10 && pixel_y < 14) || (pixel_x == 1316 && pixel_y == 10) || (pixel_x == 1322 && pixel_y >= 10 && pixel_y < 12) || (pixel_x >= 1345 && pixel_x < 1347 && pixel_y >= 10 && pixel_y < 12) || (pixel_x == 1347 && pixel_y == 10) || (pixel_x == 1359 && pixel_y == 10) || (pixel_x == 39 && pixel_y >= 11 && pixel_y < 18) || (pixel_x == 63 && pixel_y == 11) || (pixel_x == 138 && pixel_y == 11) || (pixel_x == 146 && pixel_y == 11) || (pixel_x == 217 && pixel_y >= 11 && pixel_y < 15) || (pixel_x == 232 && pixel_y >= 11 && pixel_y < 15) || (pixel_x == 263 && pixel_y >= 11 && pixel_y < 14) || (pixel_x >= 274 && pixel_x < 277 && pixel_y >= 11 && pixel_y < 13) || (pixel_x >= 309 && pixel_x < 311 && pixel_y >= 11 && pixel_y < 14) || (pixel_x >= 320 && pixel_x < 322 && pixel_y >= 11 && pixel_y < 13) || (pixel_x >= 325 && pixel_x < 327 && pixel_y >= 11 && pixel_y < 13) || (pixel_x == 363 && pixel_y >= 11 && pixel_y < 14) || (pixel_x >= 382 && pixel_x < 384 && pixel_y == 11) || (pixel_x >= 396 && pixel_x < 398 && pixel_y == 11) || (pixel_x >= 414 && pixel_x < 416 && pixel_y >= 11 && pixel_y < 13) || (pixel_x == 437 && pixel_y == 11) || (pixel_x >= 440 && pixel_x < 442 && pixel_y >= 11 && pixel_y < 13) || (pixel_x == 457 && pixel_y >= 11 && pixel_y < 15) || (pixel_x >= 502 && pixel_x < 504 && pixel_y >= 11 && pixel_y < 14) || (pixel_x >= 545 && pixel_x < 552 && pixel_y >= 11 && pixel_y < 13) || (pixel_x >= 560 && pixel_x < 567 && pixel_y >= 11 && pixel_y < 13) || (pixel_x >= 589 && pixel_x < 596 && pixel_y >= 11 && pixel_y < 13) || (pixel_x >= 634 && pixel_x < 636 && pixel_y >= 11 && pixel_y < 13) || (pixel_x == 715 && pixel_y >= 11 && pixel_y < 14) || (pixel_x >= 743 && pixel_x < 745 && pixel_y >= 11 && pixel_y < 17) || (pixel_x >= 757 && pixel_x < 759 && pixel_y >= 11 && pixel_y < 14) || (pixel_x == 800 && pixel_y >= 11 && pixel_y < 19) || (pixel_x == 918 && pixel_y >= 11 && pixel_y < 16) || (pixel_x == 926 && pixel_y >= 11 && pixel_y < 15) || (pixel_x == 964 && pixel_y >= 11 && pixel_y < 13) || (pixel_x == 993 && pixel_y >= 11 && pixel_y < 20) || (pixel_x == 1024 && pixel_y >= 11 && pixel_y < 16) || (pixel_x == 1118 && pixel_y >= 11 && pixel_y < 14) || (pixel_x == 1147 && pixel_y >= 11 && pixel_y < 22) || (pixel_x == 1172 && pixel_y >= 11 && pixel_y < 20) || (pixel_x == 1181 && pixel_y >= 11 && pixel_y < 13) || (pixel_x == 1189 && pixel_y >= 11 && pixel_y < 14) || (pixel_x == 1198 && pixel_y >= 11 && pixel_y < 16) || (pixel_x == 1203 && pixel_y >= 11 && pixel_y < 21) || (pixel_x >= 1286 && pixel_x < 1288 && pixel_y >= 11 && pixel_y < 14) || (pixel_x == 1299 && pixel_y >= 11 && pixel_y < 18) || (pixel_x == 1303 && pixel_y >= 11 && pixel_y < 17) || (pixel_x == 1311 && pixel_y >= 11 && pixel_y < 18) || (pixel_x == 1324 && pixel_y >= 11 && pixel_y < 16) || (pixel_x == 1331 && pixel_y >= 11 && pixel_y < 16) || (pixel_x == 1344 && pixel_y >= 11 && pixel_y < 15) || (pixel_x == 54 && pixel_y >= 12 && pixel_y < 15) || (pixel_x == 77 && pixel_y >= 12 && pixel_y < 16) || (pixel_x >= 86 && pixel_x < 88 && pixel_y >= 12 && pixel_y < 18) || (pixel_x == 107 && pixel_y >= 12 && pixel_y < 16) || (pixel_x == 132 && pixel_y >= 12 && pixel_y < 17) || (pixel_x == 216 && pixel_y >= 12 && pixel_y < 16) || (pixel_x == 231 && pixel_y >= 12 && pixel_y < 16) || (pixel_x == 262 && pixel_y >= 12 && pixel_y < 14) || (pixel_x >= 280 && pixel_x < 282 && pixel_y >= 12 && pixel_y < 15) || (pixel_x == 287 && pixel_y >= 12 && pixel_y < 17) || (pixel_x >= 307 && pixel_x < 309 && pixel_y == 12) || (pixel_x == 311 && pixel_y >= 12 && pixel_y < 21) || (pixel_x == 319 && pixel_y >= 12 && pixel_y < 22) || (pixel_x == 327 && pixel_y >= 12 && pixel_y < 21) || (pixel_x == 337 && pixel_y >= 12 && pixel_y < 15) || (pixel_x == 355 && pixel_y >= 12 && pixel_y < 16) || (pixel_x == 364 && pixel_y >= 12 && pixel_y < 14) || (pixel_x >= 368 && pixel_x < 370 && pixel_y >= 12 && pixel_y < 14) || (pixel_x >= 412 && pixel_x < 414 && pixel_y >= 12 && pixel_y < 14) || (pixel_x >= 421 && pixel_x < 434 && pixel_y >= 12 && pixel_y < 14) || (pixel_x == 439 && pixel_y == 12) || (pixel_x >= 442 && pixel_x < 444 && pixel_y >= 12 && pixel_y < 14) || (pixel_x == 456 && pixel_y >= 12 && pixel_y < 17) || (pixel_x == 458 && pixel_y == 12) || (pixel_x == 473 && pixel_y >= 12 && pixel_y < 15) || (pixel_x == 478 && pixel_y >= 12 && pixel_y < 16) || (pixel_x == 483 && pixel_y >= 12 && pixel_y < 20) || (pixel_x == 491 && pixel_y >= 12 && pixel_y < 20) || (pixel_x >= 500 && pixel_x < 502 && pixel_y == 12) || (pixel_x == 567 && pixel_y == 12) || (pixel_x == 666 && pixel_y >= 12 && pixel_y < 18) || (pixel_x == 683 && pixel_y >= 12 && pixel_y < 17) || (pixel_x == 714 && pixel_y >= 12 && pixel_y < 15) || (pixel_x >= 739 && pixel_x < 743 && pixel_y >= 12 && pixel_y < 14) || (pixel_x >= 759 && pixel_x < 761 && pixel_y >= 12 && pixel_y < 15) || (pixel_x == 804 && pixel_y >= 12 && pixel_y < 20) || (pixel_x == 812 && pixel_y >= 12 && pixel_y < 21) || (pixel_x == 820 && pixel_y >= 12 && pixel_y < 22) || (pixel_x == 861 && pixel_y >= 12 && pixel_y < 17) || (pixel_x == 893 && pixel_y >= 12 && pixel_y < 16) || (pixel_x == 962 && pixel_y >= 12 && pixel_y < 21) || (pixel_x == 979 && pixel_y >= 12 && pixel_y < 14) || (pixel_x == 988 && pixel_y >= 12 && pixel_y < 16) || (pixel_x == 1007 && pixel_y >= 12 && pixel_y < 20) || (pixel_x == 1009 && pixel_y == 12) || (pixel_x == 1022 && pixel_y >= 12 && pixel_y < 19) || (pixel_x == 1052 && pixel_y >= 12 && pixel_y < 20) || (pixel_x == 1054 && pixel_y == 12) || (pixel_x == 1069 && pixel_y >= 12 && pixel_y < 14) || (pixel_x == 1117 && pixel_y >= 12 && pixel_y < 17) || (pixel_x == 1148 && pixel_y >= 12 && pixel_y < 22) || (pixel_x == 1159 && pixel_y >= 12 && pixel_y < 14) || (pixel_x == 1173 && pixel_y >= 12 && pixel_y < 21) || (pixel_x == 1183 && pixel_y >= 12 && pixel_y < 18) || (pixel_x == 1202 && pixel_y >= 12 && pixel_y < 20) || (pixel_x == 1235 && pixel_y >= 12 && pixel_y < 15) || (pixel_x == 1279 && pixel_y >= 12 && pixel_y < 17) || (pixel_x >= 1312 && pixel_x < 1314 && pixel_y >= 12 && pixel_y < 17) || (pixel_x == 1332 && pixel_y >= 12 && pixel_y < 14) || (pixel_x == 1343 && pixel_y >= 12 && pixel_y < 16) || (pixel_x == 1345 && pixel_y == 12) || (pixel_x == 1356 && pixel_y >= 12 && pixel_y < 16) || (pixel_x == 1388 && pixel_y >= 12 && pixel_y < 17) || (pixel_x >= 6 && pixel_x < 8 && pixel_y >= 13 && pixel_y < 16) || (pixel_x >= 55 && pixel_x < 57 && pixel_y >= 13 && pixel_y < 16) || (pixel_x >= 69 && pixel_x < 71 && pixel_y >= 13 && pixel_y < 15) || (pixel_x >= 71 && pixel_x < 74 && pixel_y == 13) || (pixel_x == 76 && pixel_y >= 13 && pixel_y < 21) || (pixel_x >= 80 && pixel_x < 83 && pixel_y == 13) || (pixel_x >= 183 && pixel_x < 192 && pixel_y >= 13 && pixel_y < 15) || (pixel_x == 261 && pixel_y >= 13 && pixel_y < 16) || (pixel_x == 282 && pixel_y >= 13 && pixel_y < 20) || (pixel_x == 286 && pixel_y >= 13 && pixel_y < 17) || (pixel_x == 312 && pixel_y >= 13 && pixel_y < 20) || (pixel_x == 320 && pixel_y == 13) || (pixel_x == 326 && pixel_y == 13) || (pixel_x == 328 && pixel_y >= 13 && pixel_y < 19) || (pixel_x == 336 && pixel_y >= 13 && pixel_y < 19) || (pixel_x == 349 && pixel_y >= 13 && pixel_y < 16) || (pixel_x == 353 && pixel_y == 13) || (pixel_x == 356 && pixel_y >= 13 && pixel_y < 22) || (pixel_x >= 365 && pixel_x < 368 && pixel_y >= 13 && pixel_y < 15) || (pixel_x >= 410 && pixel_x < 412 && pixel_y >= 13 && pixel_y < 15) || (pixel_x == 441 && pixel_y == 13) || (pixel_x >= 444 && pixel_x < 446 && pixel_y >= 13 && pixel_y < 17) || (pixel_x >= 505 && pixel_x < 507 && pixel_y >= 13 && pixel_y < 16) || (pixel_x == 560 && pixel_y == 13) || (pixel_x >= 579 && pixel_x < 583 && pixel_y == 13) || (pixel_x == 635 && pixel_y == 13) || (pixel_x == 638 && pixel_y >= 13 && pixel_y < 18) || (pixel_x == 668 && pixel_y >= 13 && pixel_y < 18) || (pixel_x >= 710 && pixel_x < 714 && pixel_y >= 13 && pixel_y < 15) || (pixel_x == 761 && pixel_y >= 13 && pixel_y < 21) || (pixel_x == 815 && pixel_y >= 13 && pixel_y < 19) || (pixel_x == 830 && pixel_y >= 13 && pixel_y < 18) || (pixel_x == 834 && pixel_y >= 13 && pixel_y < 18) || (pixel_x == 860 && pixel_y >= 13 && pixel_y < 18) || (pixel_x == 917 && pixel_y >= 13 && pixel_y < 16) || (pixel_x == 927 && pixel_y >= 13 && pixel_y < 16) || (pixel_x == 992 && pixel_y >= 13 && pixel_y < 18) || (pixel_x == 1033 && pixel_y >= 13 && pixel_y < 15) || (pixel_x == 1116 && pixel_y >= 13 && pixel_y < 16) || (pixel_x == 1171 && pixel_y >= 13 && pixel_y < 17) || (pixel_x == 1236 && pixel_y >= 13 && pixel_y < 16) || (pixel_x == 1285 && pixel_y >= 13 && pixel_y < 18) || (pixel_x == 1295 && pixel_y >= 13 && pixel_y < 20) || (pixel_x == 1298 && pixel_y >= 13 && pixel_y < 15) || (pixel_x == 1302 && pixel_y >= 13 && pixel_y < 22) || (pixel_x == 1325 && pixel_y >= 13 && pixel_y < 18) || (pixel_x == 1330 && pixel_y >= 13 && pixel_y < 19) || (pixel_x == 1342 && pixel_y >= 13 && pixel_y < 17) || (pixel_x >= 1353 && pixel_x < 1356 && pixel_y >= 13 && pixel_y < 15) || (pixel_x >= 1389 && pixel_x < 1392 && pixel_y >= 13 && pixel_y < 15) || (pixel_x >= 1397 && pixel_x < 1402 && pixel_y >= 13 && pixel_y < 15) || (pixel_x == 1408 && pixel_y >= 13 && pixel_y < 16) || (pixel_x == 33 && pixel_y >= 14 && pixel_y < 21) || (pixel_x == 57 && pixel_y >= 14 && pixel_y < 20) || (pixel_x == 65 && pixel_y >= 14 && pixel_y < 17) || (pixel_x >= 72 && pixel_x < 74 && pixel_y == 14) || (pixel_x >= 81 && pixel_x < 84 && pixel_y == 14) || (pixel_x >= 151 && pixel_x < 157 && pixel_y >= 14 && pixel_y < 16) || (pixel_x >= 158 && pixel_x < 164 && pixel_y >= 14 && pixel_y < 16) || (pixel_x == 215 && pixel_y >= 14 && pixel_y < 18) || (pixel_x == 230 && pixel_y >= 14 && pixel_y < 18) || (pixel_x == 260 && pixel_y >= 14 && pixel_y < 17) || (pixel_x == 310 && pixel_y == 14) || (pixel_x == 348 && pixel_y >= 14 && pixel_y < 21) || (pixel_x == 357 && pixel_y >= 14 && pixel_y < 21) || (pixel_x >= 408 && pixel_x < 410 && pixel_y >= 14 && pixel_y < 17) || (pixel_x == 443 && pixel_y == 14) || (pixel_x >= 446 && pixel_x < 448 && pixel_y >= 14 && pixel_y < 16) || (pixel_x == 455 && pixel_y >= 14 && pixel_y < 17) || (pixel_x >= 470 && pixel_x < 473 && pixel_y >= 14 && pixel_y < 16) || (pixel_x == 477 && pixel_y >= 14 && pixel_y < 16) || (pixel_x >= 581 && pixel_x < 583 && pixel_y >= 14 && pixel_y < 22) || (pixel_x == 684 && pixel_y >= 14 && pixel_y < 19) || (pixel_x == 693 && pixel_y >= 14 && pixel_y < 21) || (pixel_x == 723 && pixel_y >= 14 && pixel_y < 21) || (pixel_x == 742 && pixel_y == 14) || (pixel_x == 762 && pixel_y >= 14 && pixel_y < 20) || (pixel_x == 801 && pixel_y >= 14 && pixel_y < 22) || (pixel_x == 814 && pixel_y >= 14 && pixel_y < 22) || (pixel_x == 821 && pixel_y >= 14 && pixel_y < 22) || (pixel_x == 894 && pixel_y >= 14 && pixel_y < 18) || (pixel_x >= 1025 && pixel_x < 1031 && pixel_y >= 14 && pixel_y < 16) || (pixel_x == 1115 && pixel_y == 14) || (pixel_x == 1234 && pixel_y == 14) || (pixel_x >= 1237 && pixel_x < 1240 && pixel_y >= 14 && pixel_y < 16) || (pixel_x == 1280 && pixel_y >= 14 && pixel_y < 20) || (pixel_x == 1286 && pixel_y >= 14 && pixel_y < 16) || (pixel_x == 1293 && pixel_y >= 14 && pixel_y < 22) || (pixel_x == 1300 && pixel_y >= 14 && pixel_y < 22) || (pixel_x == 1341 && pixel_y >= 14 && pixel_y < 18) || (pixel_x == 1392 && pixel_y == 14) || (pixel_x >= 1402 && pixel_x < 1404 && pixel_y >= 14 && pixel_y < 16) || (pixel_x >= 31 && pixel_x < 33 && pixel_y >= 15 && pixel_y < 17) || (pixel_x >= 35 && pixel_x < 39 && pixel_y >= 15 && pixel_y < 17) || (pixel_x >= 40 && pixel_x < 44 && pixel_y >= 15 && pixel_y < 17) || (pixel_x == 64 && pixel_y >= 15 && pixel_y < 19) || (pixel_x == 69 && pixel_y == 15) || (pixel_x >= 73 && pixel_x < 76 && pixel_y >= 15 && pixel_y < 20) || (pixel_x >= 82 && pixel_x < 85 && pixel_y == 15) || (pixel_x >= 228 && pixel_x < 230 && pixel_y >= 15 && pixel_y < 21) || (pixel_x == 236 && pixel_y >= 15 && pixel_y < 21) || (pixel_x == 259 && pixel_y >= 15 && pixel_y < 19) || (pixel_x == 281 && pixel_y >= 15 && pixel_y < 21) || (pixel_x >= 288 && pixel_x < 294 && pixel_y >= 15 && pixel_y < 17) || (pixel_x >= 296 && pixel_x < 299 && pixel_y >= 15 && pixel_y < 17) || (pixel_x == 335 && pixel_y >= 15 && pixel_y < 22) || (pixel_x == 347 && pixel_y >= 15 && pixel_y < 20) || (pixel_x >= 406 && pixel_x < 408 && pixel_y == 15) || (pixel_x == 410 && pixel_y >= 15 && pixel_y < 18) || (pixel_x == 448 && pixel_y == 15) || (pixel_x == 469 && pixel_y == 15) || (pixel_x == 476 && pixel_y >= 15 && pixel_y < 17) || (pixel_x == 482 && pixel_y >= 15 && pixel_y < 22) || (pixel_x == 492 && pixel_y >= 15 && pixel_y < 22) || (pixel_x == 507 && pixel_y >= 15 && pixel_y < 20) || (pixel_x == 536 && pixel_y >= 15 && pixel_y < 20) || (pixel_x == 639 && pixel_y >= 15 && pixel_y < 19) || (pixel_x == 667 && pixel_y >= 15 && pixel_y < 18) || (pixel_x == 745 && pixel_y >= 15 && pixel_y < 20) || (pixel_x == 760 && pixel_y == 15) || (pixel_x == 829 && pixel_y >= 15 && pixel_y < 20) || (pixel_x == 835 && pixel_y >= 15 && pixel_y < 20) || (pixel_x == 859 && pixel_y >= 15 && pixel_y < 22) || (pixel_x == 895 && pixel_y >= 15 && pixel_y < 19) || (pixel_x == 916 && pixel_y == 15) || (pixel_x == 928 && pixel_y == 15) || (pixel_x == 961 && pixel_y >= 15 && pixel_y < 18) || (pixel_x == 1118 && pixel_y >= 15 && pixel_y < 19) || (pixel_x >= 1240 && pixel_x < 1242 && pixel_y >= 15 && pixel_y < 18) || (pixel_x == 1284 && pixel_y >= 15 && pixel_y < 21) || (pixel_x == 1314 && pixel_y >= 15 && pixel_y < 19) || (pixel_x == 1326 && pixel_y >= 15 && pixel_y < 20) || (pixel_x >= 1357 && pixel_x < 1359 && pixel_y >= 15 && pixel_y < 25) || (pixel_x == 1387 && pixel_y >= 15 && pixel_y < 26) || (pixel_x == 1389 && pixel_y == 15) || (pixel_x >= 1396 && pixel_x < 1398 && pixel_y == 15) || (pixel_x == 1401 && pixel_y == 15) || (pixel_x >= 1404 && pixel_x < 1408 && pixel_y >= 15 && pixel_y < 17) || (pixel_x == 7 && pixel_y == 16) || (pixel_x == 56 && pixel_y >= 16 && pixel_y < 21) || (pixel_x == 67 && pixel_y >= 16 && pixel_y < 19) || (pixel_x >= 83 && pixel_x < 86 && pixel_y >= 16 && pixel_y < 18) || (pixel_x == 156 && pixel_y == 16) || (pixel_x == 158 && pixel_y == 16) || (pixel_x == 214 && pixel_y >= 16 && pixel_y < 20) || (pixel_x == 258 && pixel_y >= 16 && pixel_y < 22) || (pixel_x == 313 && pixel_y == 16) || (pixel_x == 411 && pixel_y >= 16 && pixel_y < 18) || (pixel_x == 443 && pixel_y >= 16 && pixel_y < 18) || (pixel_x == 446 && pixel_y == 16) || (pixel_x == 470 && pixel_y == 16) || (pixel_x >= 485 && pixel_x < 490 && pixel_y >= 16 && pixel_y < 18) || (pixel_x == 506 && pixel_y >= 16 && pixel_y < 21) || (pixel_x == 514 && pixel_y >= 16 && pixel_y < 21) || (pixel_x == 574 && pixel_y >= 16 && pixel_y < 21) || (pixel_x == 640 && pixel_y >= 16 && pixel_y < 20) || (pixel_x == 685 && pixel_y >= 16 && pixel_y < 20) || (pixel_x == 701 && pixel_y >= 16 && pixel_y < 21) || (pixel_x == 731 && pixel_y >= 16 && pixel_y < 21) || (pixel_x == 763 && pixel_y >= 16 && pixel_y < 18) || (pixel_x == 803 && pixel_y >= 16 && pixel_y < 22) || (pixel_x == 836 && pixel_y >= 16 && pixel_y < 22) || (pixel_x == 1119 && pixel_y >= 16 && pixel_y < 20) || (pixel_x == 1239 && pixel_y == 16) || (pixel_x == 1242 && pixel_y >= 16 && pixel_y < 21) || (pixel_x == 1281 && pixel_y >= 16 && pixel_y < 22) || (pixel_x == 1310 && pixel_y >= 16 && pixel_y < 19) || (pixel_x == 1329 && pixel_y >= 16 && pixel_y < 21) || (pixel_x == 1340 && pixel_y >= 16 && pixel_y < 19) || (pixel_x == 1386 && pixel_y >= 16 && pixel_y < 22) || (pixel_x == 1396 && pixel_y == 16) || (pixel_x == 1403 && pixel_y == 16) || (pixel_x == 38 && pixel_y >= 17 && pixel_y < 22) || (pixel_x == 63 && pixel_y >= 17 && pixel_y < 20) || (pixel_x == 213 && pixel_y >= 17 && pixel_y < 21) || (pixel_x == 334 && pixel_y >= 17 && pixel_y < 22) || (pixel_x == 358 && pixel_y >= 17 && pixel_y < 19) || (pixel_x >= 412 && pixel_x < 414 && pixel_y >= 17 && pixel_y < 19) || (pixel_x >= 421 && pixel_x < 434 && pixel_y == 17) || (pixel_x >= 441 && pixel_x < 443 && pixel_y >= 17 && pixel_y < 19) || (pixel_x == 444 && pixel_y == 17) || (pixel_x == 467 && pixel_y >= 17 && pixel_y < 20) || (pixel_x == 641 && pixel_y >= 17 && pixel_y < 21) || (pixel_x == 744 && pixel_y == 17) || (pixel_x == 746 && pixel_y >= 17 && pixel_y < 21) || (pixel_x >= 791 && pixel_x < 793 && pixel_y >= 17 && pixel_y < 20) || (pixel_x == 802 && pixel_y >= 17 && pixel_y < 22) || (pixel_x == 828 && pixel_y >= 17 && pixel_y < 22) || (pixel_x == 858 && pixel_y >= 17 && pixel_y < 22) || (pixel_x == 896 && pixel_y >= 17 && pixel_y < 21) || (pixel_x == 970 && pixel_y >= 17 && pixel_y < 20) || (pixel_x == 1015 && pixel_y >= 17 && pixel_y < 20) || (pixel_x == 1024 && pixel_y >= 17 && pixel_y < 21) || (pixel_x == 1060 && pixel_y >= 17 && pixel_y < 20) || (pixel_x == 1120 && pixel_y >= 17 && pixel_y < 21) || (pixel_x == 1181 && pixel_y >= 17 && pixel_y < 21) || (pixel_x == 1210 && pixel_y >= 17 && pixel_y < 20) || (pixel_x == 1270 && pixel_y >= 17 && pixel_y < 20) || (pixel_x == 1294 && pixel_y >= 17 && pixel_y < 22) || (pixel_x == 1301 && pixel_y >= 17 && pixel_y < 22) || (pixel_x == 1309 && pixel_y >= 17 && pixel_y < 21) || (pixel_x == 1313 && pixel_y == 17) || (pixel_x == 1315 && pixel_y >= 17 && pixel_y < 20) || (pixel_x == 1327 && pixel_y >= 17 && pixel_y < 25) || (pixel_x == 1339 && pixel_y >= 17 && pixel_y < 22) || (pixel_x == 1359 && pixel_y >= 17 && pixel_y < 19) || (pixel_x == 32 && pixel_y >= 18 && pixel_y < 22) || (pixel_x >= 84 && pixel_x < 87 && pixel_y >= 18 && pixel_y < 21) || (pixel_x == 110 && pixel_y >= 18 && pixel_y < 23) || (pixel_x == 129 && pixel_y >= 18 && pixel_y < 23) || (pixel_x == 172 && pixel_y >= 18 && pixel_y < 26) || (pixel_x == 257 && pixel_y >= 18 && pixel_y < 22) || (pixel_x == 280 && pixel_y >= 18 && pixel_y < 22) || (pixel_x == 310 && pixel_y >= 18 && pixel_y < 22) || (pixel_x == 326 && pixel_y >= 18 && pixel_y < 21) || (pixel_x == 349 && pixel_y >= 18 && pixel_y < 22) || (pixel_x == 370 && pixel_y >= 18 && pixel_y < 21) || (pixel_x == 397 && pixel_y >= 18 && pixel_y < 26) || (pixel_x >= 414 && pixel_x < 416 && pixel_y >= 18 && pixel_y < 20) || (pixel_x >= 439 && pixel_x < 441 && pixel_y >= 18 && pixel_y < 20) || (pixel_x == 493 && pixel_y >= 18 && pixel_y < 22) || (pixel_x == 505 && pixel_y >= 18 && pixel_y < 21) || (pixel_x == 515 && pixel_y >= 18 && pixel_y < 21) || (pixel_x == 535 && pixel_y >= 18 && pixel_y < 21) || (pixel_x == 575 && pixel_y >= 18 && pixel_y < 21) || (pixel_x == 694 && pixel_y >= 18 && pixel_y < 22) || (pixel_x == 724 && pixel_y >= 18 && pixel_y < 22) || (pixel_x == 747 && pixel_y >= 18 && pixel_y < 22) || (pixel_x == 837 && pixel_y >= 18 && pixel_y < 22) || (pixel_x == 857 && pixel_y >= 18 && pixel_y < 22) || (pixel_x == 969 && pixel_y >= 18 && pixel_y < 21) || (pixel_x == 985 && pixel_y >= 18 && pixel_y < 21) || (pixel_x == 995 && pixel_y >= 18 && pixel_y < 21) || (pixel_x == 1014 && pixel_y >= 18 && pixel_y < 21) || (pixel_x == 1121 && pixel_y >= 18 && pixel_y < 22) || (pixel_x == 1174 && pixel_y >= 18 && pixel_y < 22) || (pixel_x == 1195 && pixel_y >= 18 && pixel_y < 21) || (pixel_x == 1241 && pixel_y >= 18 && pixel_y < 22) || (pixel_x == 1269 && pixel_y >= 18 && pixel_y < 21) || (pixel_x >= 1282 && pixel_x < 1284 && pixel_y >= 18 && pixel_y < 22) || (pixel_x == 1308 && pixel_y >= 18 && pixel_y < 22) || (pixel_x == 1316 && pixel_y >= 18 && pixel_y < 22) || (pixel_x == 1328 && pixel_y >= 18 && pixel_y < 23) || (pixel_x == 1338 && pixel_y >= 18 && pixel_y < 22) || (pixel_x >= 6 && pixel_x < 9 && pixel_y >= 19 && pixel_y < 22) || (pixel_x == 37 && pixel_y >= 19 && pixel_y < 22) || (pixel_x >= 47 && pixel_x < 49 && pixel_y >= 19 && pixel_y < 21) || (pixel_x >= 54 && pixel_x < 56 && pixel_y >= 19 && pixel_y < 21) || (pixel_x == 62 && pixel_y >= 19 && pixel_y < 22) || (pixel_x == 69 && pixel_y >= 19 && pixel_y < 22) || (pixel_x == 72 && pixel_y >= 19 && pixel_y < 22) || (pixel_x == 77 && pixel_y >= 19 && pixel_y < 22) || (pixel_x == 87 && pixel_y >= 19 && pixel_y < 22) || (pixel_x == 171 && pixel_y >= 19 && pixel_y < 22) || (pixel_x == 173 && pixel_y >= 19 && pixel_y < 25) || (pixel_x >= 201 && pixel_x < 204 && pixel_y >= 19 && pixel_y < 22) || (pixel_x == 212 && pixel_y >= 19 && pixel_y < 23) || (pixel_x == 235 && pixel_y >= 19 && pixel_y < 22) || (pixel_x == 302 && pixel_y >= 19 && pixel_y < 22) || (pixel_x == 309 && pixel_y >= 19 && pixel_y < 22) || (pixel_x == 320 && pixel_y >= 19 && pixel_y < 22) || (pixel_x == 325 && pixel_y >= 19 && pixel_y < 22) || (pixel_x == 355 && pixel_y >= 19 && pixel_y < 22) || (pixel_x == 369 && pixel_y >= 19 && pixel_y < 22) || (pixel_x >= 381 && pixel_x < 384 && pixel_y >= 19 && pixel_y < 22) || (pixel_x == 396 && pixel_y >= 19 && pixel_y < 22) || (pixel_x == 398 && pixel_y >= 19 && pixel_y < 25) || (pixel_x >= 416 && pixel_x < 418 && pixel_y >= 19 && pixel_y < 21) || (pixel_x >= 437 && pixel_x < 439 && pixel_y >= 19 && pixel_y < 21) || (pixel_x >= 455 && pixel_x < 457 && pixel_y >= 19 && pixel_y < 22) || (pixel_x == 468 && pixel_y >= 19 && pixel_y < 21) || (pixel_x == 481 && pixel_y >= 19 && pixel_y < 22) || (pixel_x == 504 && pixel_y >= 19 && pixel_y < 22) || (pixel_x == 516 && pixel_y >= 19 && pixel_y < 22) || (pixel_x == 534 && pixel_y >= 19 && pixel_y < 22) || (pixel_x == 576 && pixel_y >= 19 && pixel_y < 22) || (pixel_x >= 623 && pixel_x < 625 && pixel_y >= 19 && pixel_y < 21) || (pixel_x == 625 && pixel_y == 19) || (pixel_x == 642 && pixel_y >= 19 && pixel_y < 22) || (pixel_x == 700 && pixel_y >= 19 && pixel_y < 22) || (pixel_x == 730 && pixel_y >= 19 && pixel_y < 22) || (pixel_x == 752 && pixel_y >= 19 && pixel_y < 22) || (pixel_x == 760 && pixel_y >= 19 && pixel_y < 22) || (pixel_x == 784 && pixel_y >= 19 && pixel_y < 22) || (pixel_x == 790 && pixel_y >= 19 && pixel_y < 22) || (pixel_x == 827 && pixel_y >= 19 && pixel_y < 22) || (pixel_x == 897 && pixel_y >= 19 && pixel_y < 22) || (pixel_x == 964 && pixel_y >= 19 && pixel_y < 22) || (pixel_x == 968 && pixel_y >= 19 && pixel_y < 21) || (pixel_x == 984 && pixel_y >= 19 && pixel_y < 22) || (pixel_x == 996 && pixel_y >= 19 && pixel_y < 22) || (pixel_x == 1009 && pixel_y >= 19 && pixel_y < 22) || (pixel_x == 1013 && pixel_y >= 19 && pixel_y < 22) || (pixel_x == 1025 && pixel_y >= 19 && pixel_y < 22) || (pixel_x == 1032 && pixel_y >= 19 && pixel_y < 21) || (pixel_x == 1054 && pixel_y >= 19 && pixel_y < 22) || (pixel_x >= 1058 && pixel_x < 1060 && pixel_y >= 19 && pixel_y < 21) || (pixel_x == 1180 && pixel_y >= 19 && pixel_y < 22) || (pixel_x == 1194 && pixel_y >= 19 && pixel_y < 22) || (pixel_x == 1196 && pixel_y == 19) || (pixel_x == 1204 && pixel_y >= 19 && pixel_y < 22) || (pixel_x >= 1208 && pixel_x < 1210 && pixel_y >= 19 && pixel_y < 21) || (pixel_x == 1232 && pixel_y >= 19 && pixel_y < 21) || (pixel_x == 1240 && pixel_y >= 19 && pixel_y < 22) || (pixel_x == 1252 && pixel_y >= 19 && pixel_y < 22) || (pixel_x == 1264 && pixel_y >= 19 && pixel_y < 22) || (pixel_x == 1268 && pixel_y >= 19 && pixel_y < 22) || (pixel_x == 1317 && pixel_y >= 19 && pixel_y < 22) || (pixel_x == 1337 && pixel_y >= 19 && pixel_y < 22) || (pixel_x >= 49 && pixel_x < 52 && pixel_y >= 20 && pixel_y < 22) || (pixel_x == 61 && pixel_y >= 20 && pixel_y < 23) || (pixel_x >= 70 && pixel_x < 72 && pixel_y >= 20 && pixel_y < 22) || (pixel_x == 73 && pixel_y == 20) || (pixel_x >= 78 && pixel_x < 80 && pixel_y >= 20 && pixel_y < 22) || (pixel_x >= 82 && pixel_x < 84 && pixel_y >= 20 && pixel_y < 22) || (pixel_x == 88 && pixel_y >= 20 && pixel_y < 22) || (pixel_x == 111 && pixel_y >= 20 && pixel_y < 24) || (pixel_x == 128 && pixel_y >= 20 && pixel_y < 24) || (pixel_x == 170 && pixel_y == 20) || (pixel_x == 174 && pixel_y >= 20 && pixel_y < 23) || (pixel_x >= 230 && pixel_x < 232 && pixel_y >= 20 && pixel_y < 22) || (pixel_x >= 233 && pixel_x < 235 && pixel_y >= 20 && pixel_y < 22) || (pixel_x >= 242 && pixel_x < 247 && pixel_y >= 20 && pixel_y < 22) || (pixel_x >= 249 && pixel_x < 254 && pixel_y >= 20 && pixel_y < 22) || (pixel_x >= 259 && pixel_x < 268 && pixel_y >= 20 && pixel_y < 22) || (pixel_x >= 272 && pixel_x < 275 && pixel_y >= 20 && pixel_y < 22) || (pixel_x >= 278 && pixel_x < 280 && pixel_y >= 20 && pixel_y < 22) || (pixel_x >= 303 && pixel_x < 309 && pixel_y >= 20 && pixel_y < 22) || (pixel_x >= 321 && pixel_x < 323 && pixel_y >= 20 && pixel_y < 22) || (pixel_x == 324 && pixel_y >= 20 && pixel_y < 22) || (pixel_x >= 350 && pixel_x < 352 && pixel_y >= 20 && pixel_y < 22) || (pixel_x >= 353 && pixel_x < 355 && pixel_y >= 20 && pixel_y < 22) || (pixel_x >= 362 && pixel_x < 365 && pixel_y >= 20 && pixel_y < 22) || (pixel_x >= 367 && pixel_x < 369 && pixel_y >= 20 && pixel_y < 22) || (pixel_x == 395 && pixel_y == 20) || (pixel_x == 399 && pixel_y >= 20 && pixel_y < 23) || (pixel_x == 418 && pixel_y >= 20 && pixel_y < 22) || (pixel_x == 436 && pixel_y >= 20 && pixel_y < 22) || (pixel_x == 457 && pixel_y >= 20 && pixel_y < 22) || (pixel_x == 469 && pixel_y >= 20 && pixel_y < 22) || (pixel_x == 475 && pixel_y >= 20 && pixel_y < 22) || (pixel_x >= 500 && pixel_x < 504 && pixel_y >= 20 && pixel_y < 22) || (pixel_x >= 517 && pixel_x < 519 && pixel_y >= 20 && pixel_y < 22) || (pixel_x >= 521 && pixel_x < 523 && pixel_y >= 20 && pixel_y < 22) || (pixel_x >= 529 && pixel_x < 534 && pixel_y >= 20 && pixel_y < 22) || (pixel_x >= 545 && pixel_x < 553 && pixel_y >= 20 && pixel_y < 22) || (pixel_x >= 577 && pixel_x < 579 && pixel_y >= 20 && pixel_y < 22) || (pixel_x >= 602 && pixel_x < 606 && pixel_y >= 20 && pixel_y < 22) || (pixel_x >= 609 && pixel_x < 613 && pixel_y >= 20 && pixel_y < 22) || (pixel_x >= 616 && pixel_x < 620 && pixel_y == 20) || (pixel_x == 622 && pixel_y >= 20 && pixel_y < 22) || (pixel_x == 643 && pixel_y >= 20 && pixel_y < 22) || (pixel_x >= 650 && pixel_x < 658 && pixel_y >= 20 && pixel_y < 22) || (pixel_x >= 695 && pixel_x < 697 && pixel_y >= 20 && pixel_y < 22) || (pixel_x == 699 && pixel_y >= 20 && pixel_y < 22) || (pixel_x >= 725 && pixel_x < 727 && pixel_y >= 20 && pixel_y < 22) || (pixel_x == 729 && pixel_y >= 20 && pixel_y < 26) || (pixel_x == 748 && pixel_y >= 20 && pixel_y < 22) || (pixel_x >= 753 && pixel_x < 756 && pixel_y >= 20 && pixel_y < 22) || (pixel_x >= 758 && pixel_x < 760 && pixel_y >= 20 && pixel_y < 22) || (pixel_x == 783 && pixel_y == 20) || (pixel_x >= 785 && pixel_x < 787 && pixel_y >= 20 && pixel_y < 22) || (pixel_x >= 788 && pixel_x < 790 && pixel_y >= 20 && pixel_y < 22) || (pixel_x == 791 && pixel_y == 20) || (pixel_x == 838 && pixel_y >= 20 && pixel_y < 22) || (pixel_x >= 860 && pixel_x < 869 && pixel_y >= 20 && pixel_y < 22) || (pixel_x == 898 && pixel_y >= 20 && pixel_y < 23) || (pixel_x >= 965 && pixel_x < 968 && pixel_y >= 20 && pixel_y < 22) || (pixel_x >= 979 && pixel_x < 984 && pixel_y >= 20 && pixel_y < 22) || (pixel_x >= 997 && pixel_x < 1003 && pixel_y >= 20 && pixel_y < 22) || (pixel_x == 1003 && pixel_y == 20) || (pixel_x >= 1010 && pixel_x < 1013 && pixel_y >= 20 && pixel_y < 22) || (pixel_x >= 1026 && pixel_x < 1032 && pixel_y >= 20 && pixel_y < 22) || (pixel_x >= 1055 && pixel_x < 1058 && pixel_y >= 20 && pixel_y < 22) || (pixel_x >= 1088 && pixel_x < 1092 && pixel_y >= 20 && pixel_y < 22) || (pixel_x == 1122 && pixel_y >= 20 && pixel_y < 22) || (pixel_x >= 1133 && pixel_x < 1137 && pixel_y >= 20 && pixel_y < 22) || (pixel_x >= 1175 && pixel_x < 1180 && pixel_y >= 20 && pixel_y < 22) || (pixel_x >= 1189 && pixel_x < 1194 && pixel_y >= 20 && pixel_y < 22) || (pixel_x >= 1205 && pixel_x < 1208 && pixel_y >= 20 && pixel_y < 22) || (pixel_x >= 1233 && pixel_x < 1240 && pixel_y >= 20 && pixel_y < 22) || (pixel_x == 1251 && pixel_y == 20) || (pixel_x >= 1253 && pixel_x < 1258 && pixel_y >= 20 && pixel_y < 22) || (pixel_x == 1263 && pixel_y == 20) || (pixel_x >= 1265 && pixel_x < 1268 && pixel_y >= 20 && pixel_y < 22) || (pixel_x == 1307 && pixel_y >= 20 && pixel_y < 22) || (pixel_x == 1318 && pixel_y >= 20 && pixel_y < 22) || (pixel_x >= 1340 && pixel_x < 1348 && pixel_y >= 20 && pixel_y < 22) || (pixel_x == 1388 && pixel_y >= 20 && pixel_y < 24) || (pixel_x == 48 && pixel_y == 21) || (pixel_x == 54 && pixel_y == 21) || (pixel_x >= 80 && pixel_x < 82 && pixel_y == 21) || (pixel_x == 89 && pixel_y == 21) || (pixel_x == 211 && pixel_y >= 21 && pixel_y < 23) || (pixel_x == 229 && pixel_y == 21) || (pixel_x == 232 && pixel_y >= 21 && pixel_y < 23) || (pixel_x >= 275 && pixel_x < 278 && pixel_y == 21) || (pixel_x == 323 && pixel_y >= 21 && pixel_y < 23) || (pixel_x == 352 && pixel_y >= 21 && pixel_y < 23) || (pixel_x >= 365 && pixel_x < 367 && pixel_y >= 21 && pixel_y < 23) || (pixel_x >= 470 && pixel_x < 475 && pixel_y == 21) || (pixel_x == 494 && pixel_y == 21) || (pixel_x >= 519 && pixel_x < 521 && pixel_y == 21) || (pixel_x >= 579 && pixel_x < 581 && pixel_y >= 21 && pixel_y < 23) || (pixel_x >= 617 && pixel_x < 622 && pixel_y == 21) || (pixel_x == 623 && pixel_y == 21) || (pixel_x == 644 && pixel_y == 21) || (pixel_x >= 697 && pixel_x < 699 && pixel_y == 21) || (pixel_x >= 727 && pixel_x < 729 && pixel_y >= 21 && pixel_y < 23) || (pixel_x == 749 && pixel_y == 21) || (pixel_x >= 756 && pixel_x < 758 && pixel_y >= 21 && pixel_y < 23) || (pixel_x == 787 && pixel_y >= 21 && pixel_y < 23) || (pixel_x == 826 && pixel_y == 21) || (pixel_x == 973 && pixel_y == 21) || (pixel_x == 1058 && pixel_y == 21) || (pixel_x == 1123 && pixel_y == 21) || (pixel_x == 1208 && pixel_y == 21) || (pixel_x == 1306 && pixel_y == 21) || (pixel_x == 60 && pixel_y == 22) || (pixel_x == 80 && pixel_y == 22) || (pixel_x == 112 && pixel_y >= 22 && pixel_y < 25) || (pixel_x == 127 && pixel_y >= 22 && pixel_y < 25) || (pixel_x == 276 && pixel_y == 22) || (pixel_x >= 306 && pixel_x < 308 && pixel_y == 22) || (pixel_x == 322 && pixel_y == 22) || (pixel_x == 353 && pixel_y == 22) || (pixel_x == 472 && pixel_y == 22) || (pixel_x == 519 && pixel_y == 22) || (pixel_x >= 620 && pixel_x < 622 && pixel_y == 22) || (pixel_x == 697 && pixel_y == 22) || (pixel_x >= 931 && pixel_x < 944 && pixel_y >= 22 && pixel_y < 24) || (pixel_x >= 113 && pixel_x < 115 && pixel_y >= 23 && pixel_y < 25) || (pixel_x >= 125 && pixel_x < 127 && pixel_y >= 23 && pixel_y < 25) || (pixel_x == 728 && pixel_y >= 23 && pixel_y < 25) || (pixel_x == 1326 && pixel_y >= 23 && pixel_y < 26) || (pixel_x == 1386 && pixel_y >= 23 && pixel_y < 26) || (pixel_x >= 115 && pixel_x < 117 && pixel_y >= 24 && pixel_y < 26) || (pixel_x >= 123 && pixel_x < 125 && pixel_y >= 24 && pixel_y < 26) || (pixel_x == 730 && pixel_y >= 24 && pixel_y < 26) || (pixel_x == 908 && pixel_y >= 24 && pixel_y < 27) || (pixel_x == 1060 && pixel_y >= 24 && pixel_y < 27) || (pixel_x == 1103 && pixel_y >= 24 && pixel_y < 27) || (pixel_x == 1325 && pixel_y >= 24 && pixel_y < 27) || (pixel_x == 1359 && pixel_y >= 24 && pixel_y < 26) || (pixel_x == 1385 && pixel_y >= 24 && pixel_y < 26) || (pixel_x == 114 && pixel_y == 25) || (pixel_x == 117 && pixel_y == 25) || (pixel_x == 122 && pixel_y == 25) || (pixel_x == 125 && pixel_y == 25) || (pixel_x == 171 && pixel_y >= 25 && pixel_y < 27) || (pixel_x == 396 && pixel_y >= 25 && pixel_y < 27) || (pixel_x >= 731 && pixel_x < 735 && pixel_y >= 25 && pixel_y < 27) || (pixel_x >= 877 && pixel_x < 884 && pixel_y >= 25 && pixel_y < 27) || (pixel_x >= 901 && pixel_x < 908 && pixel_y >= 25 && pixel_y < 27) || (pixel_x >= 1052 && pixel_x < 1055 && pixel_y >= 25 && pixel_y < 27) || (pixel_x >= 1058 && pixel_x < 1060 && pixel_y >= 25 && pixel_y < 27) || (pixel_x == 1061 && pixel_y == 25) || (pixel_x == 1102 && pixel_y >= 25 && pixel_y < 27) || (pixel_x == 1104 && pixel_y == 25) || (pixel_x == 1324 && pixel_y >= 25 && pixel_y < 27) || (pixel_x == 1358 && pixel_y == 25) || (pixel_x >= 1360 && pixel_x < 1364 && pixel_y == 25) || (pixel_x >= 1382 && pixel_x < 1384 && pixel_y >= 25 && pixel_y < 27) || (pixel_x == 1384 && pixel_y == 25) || (pixel_x == 170 && pixel_y == 26) || (pixel_x == 395 && pixel_y == 26) || (pixel_x >= 875 && pixel_x < 877 && pixel_y == 26) || (pixel_x >= 1055 && pixel_x < 1058 && pixel_y >= 26 && pixel_y < 28) || (pixel_x >= 1097 && pixel_x < 1102 && pixel_y == 26) || (pixel_x >= 1321 && pixel_x < 1324 && pixel_y >= 26 && pixel_y < 28) || (pixel_x >= 1361 && pixel_x < 1363 && pixel_y == 26) || (pixel_x >= 1098 && pixel_x < 1102 && pixel_y == 27))
    hit = 1;
else hit = 0;

endmodule
