module ASCIIRenderer (
  input [10:0] x, y,
  input [7:0] ascii,
  output reg hit
);

reg [10:0] pixel_x, pixel_y;

always @ (ascii or x or y)
begin
  pixel_x = (ascii - 33) + x;
  pixel_y = y;
end

always @ (*)
if((pixel_x == 2 && pixel_y >= 1 && pixel_y < 5) || (pixel_x == 7 && pixel_y == 1) || (pixel_x == 9 && pixel_y == 1) || (pixel_x >= 18 && pixel_x < 20 && pixel_y == 1) || (pixel_x >= 22 && pixel_x < 24 && pixel_y == 1) || (pixel_x >= 28 && pixel_x < 30 && pixel_y == 1) || (pixel_x == 34 && pixel_y >= 1 && pixel_y < 3) || (pixel_x >= 40 && pixel_x < 42 && pixel_y == 1) || (pixel_x >= 44 && pixel_x < 46 && pixel_y == 1) || (pixel_x == 50 && pixel_y >= 1 && pixel_y < 5) || (pixel_x == 79 && pixel_y == 1) || (pixel_x >= 81 && pixel_x < 84 && pixel_y == 1) || (pixel_x >= 87 && pixel_x < 89 && pixel_y >= 1 && pixel_y < 3) || (pixel_x >= 92 && pixel_x < 95 && pixel_y == 1) || (pixel_x >= 97 && pixel_x < 100 && pixel_y == 1) || (pixel_x >= 104 && pixel_x < 106 && pixel_y >= 1 && pixel_y < 3) || (pixel_x >= 108 && pixel_x < 111 && pixel_y == 1) || (pixel_x >= 114 && pixel_x < 117 && pixel_y == 1) || (pixel_x >= 119 && pixel_x < 123 && pixel_y == 1) || (pixel_x >= 124 && pixel_x < 127 && pixel_y == 1) || (pixel_x >= 129 && pixel_x < 132 && pixel_y == 1) || (pixel_x >= 162 && pixel_x < 165 && pixel_y == 1) || (pixel_x == 167 && pixel_y == 1) || (pixel_x == 169 && pixel_y == 1) || (pixel_x >= 173 && pixel_x < 175 && pixel_y >= 1 && pixel_y < 4) || (pixel_x >= 177 && pixel_x < 180 && pixel_y == 1) || (pixel_x >= 184 && pixel_x < 186 && pixel_y == 1) || (pixel_x >= 188 && pixel_x < 191 && pixel_y == 1) || (pixel_x >= 194 && pixel_x < 197 && pixel_y == 1) || (pixel_x >= 199 && pixel_x < 202 && pixel_y == 1) || (pixel_x >= 205 && pixel_x < 208 && pixel_y == 1) || (pixel_x == 209 && pixel_y >= 1 && pixel_y < 8) || (pixel_x == 213 && pixel_y >= 1 && pixel_y < 7) || (pixel_x >= 215 && pixel_x < 218 && pixel_y == 1) || (pixel_x >= 221 && pixel_x < 224 && pixel_y == 1) || (pixel_x == 225 && pixel_y >= 1 && pixel_y < 7) || (pixel_x == 228 && pixel_y >= 1 && pixel_y < 3) || (pixel_x == 231 && pixel_y >= 1 && pixel_y < 8) || (pixel_x == 236 && pixel_y >= 1 && pixel_y < 7) || (pixel_x == 241 && pixel_y >= 1 && pixel_y < 7) || (pixel_x == 245 && pixel_y >= 1 && pixel_y < 5) || (pixel_x >= 247 && pixel_x < 250 && pixel_y == 1) || (pixel_x >= 252 && pixel_x < 256 && pixel_y == 1) || (pixel_x >= 258 && pixel_x < 261 && pixel_y == 1) || (pixel_x >= 263 && pixel_x < 266 && pixel_y == 1) || (pixel_x >= 269 && pixel_x < 272 && pixel_y == 1) || (pixel_x >= 273 && pixel_x < 278 && pixel_y == 1) || (pixel_x == 279 && pixel_y >= 1 && pixel_y < 8) || (pixel_x == 282 && pixel_y >= 1 && pixel_y < 7) || (pixel_x == 284 && pixel_y >= 1 && pixel_y < 3) || (pixel_x >= 288 && pixel_x < 290 && pixel_y == 1) || (pixel_x == 291 && pixel_y >= 1 && pixel_y < 4) || (pixel_x == 295 && pixel_y >= 1 && pixel_y < 3) || (pixel_x == 298 && pixel_y >= 1 && pixel_y < 3) || (pixel_x == 300 && pixel_y == 1) || (pixel_x == 304 && pixel_y == 1) || (pixel_x >= 306 && pixel_x < 310 && pixel_y == 1) || (pixel_x == 312 && pixel_y >= 1 && pixel_y < 10) || (pixel_x == 314 && pixel_y == 1) || (pixel_x == 316 && pixel_y == 1) || (pixel_x == 322 && pixel_y == 1) || (pixel_x == 324 && pixel_y >= 1 && pixel_y < 10) || (pixel_x == 339 && pixel_y == 1) || (pixel_x == 348 && pixel_y >= 1 && pixel_y < 3) || (pixel_x == 362 && pixel_y >= 1 && pixel_y < 8) || (pixel_x >= 372 && pixel_x < 374 && pixel_y == 1) || (pixel_x == 381 && pixel_y >= 1 && pixel_y < 7) || (pixel_x == 394 && pixel_y == 1) || (pixel_x == 397 && pixel_y >= 1 && pixel_y < 8) || (pixel_x == 403 && pixel_y >= 1 && pixel_y < 8) || (pixel_x >= 484 && pixel_x < 486 && pixel_y == 1) || (pixel_x == 489 && pixel_y >= 1 && pixel_y < 8) || (pixel_x == 494 && pixel_y == 1) || (pixel_x == 12 && pixel_y >= 2 && pixel_y < 6) || (pixel_x == 14 && pixel_y >= 2 && pixel_y < 6) || (pixel_x == 17 && pixel_y >= 2 && pixel_y < 4) || (pixel_x == 21 && pixel_y >= 2 && pixel_y < 4) || (pixel_x == 25 && pixel_y == 2) || (pixel_x == 27 && pixel_y == 2) || (pixel_x == 29 && pixel_y >= 2 && pixel_y < 4) || (pixel_x == 39 && pixel_y >= 2 && pixel_y < 4) || (pixel_x >= 45 && pixel_x < 47 && pixel_y == 2) || (pixel_x == 49 && pixel_y >= 2 && pixel_y < 4) || (pixel_x == 51 && pixel_y >= 2 && pixel_y < 4) || (pixel_x == 78 && pixel_y >= 2 && pixel_y < 4) || (pixel_x == 81 && pixel_y >= 2 && pixel_y < 4) || (pixel_x == 84 && pixel_y >= 2 && pixel_y < 7) || (pixel_x == 95 && pixel_y == 2) || (pixel_x == 100 && pixel_y == 2) || (pixel_x == 108 && pixel_y >= 2 && pixel_y < 4) || (pixel_x == 113 && pixel_y >= 2 && pixel_y < 7) || (pixel_x >= 121 && pixel_x < 123 && pixel_y == 2) || (pixel_x == 124 && pixel_y >= 2 && pixel_y < 4) || (pixel_x == 127 && pixel_y == 2) || (pixel_x == 129 && pixel_y >= 2 && pixel_y < 5) || (pixel_x == 132 && pixel_y >= 2 && pixel_y < 7) || (pixel_x == 164 && pixel_y >= 2 && pixel_y < 4) || (pixel_x == 166 && pixel_y >= 2 && pixel_y < 7) || (pixel_x == 170 && pixel_y == 2) || (pixel_x == 177 && pixel_y >= 2 && pixel_y < 8) || (pixel_x == 180 && pixel_y >= 2 && pixel_y < 8) || (pixel_x == 183 && pixel_y >= 2 && pixel_y < 4) || (pixel_x == 188 && pixel_y >= 2 && pixel_y < 8) || (pixel_x == 191 && pixel_y >= 2 && pixel_y < 7) || (pixel_x == 194 && pixel_y >= 2 && pixel_y < 8) || (pixel_x == 199 && pixel_y >= 2 && pixel_y < 8) || (pixel_x == 204 && pixel_y >= 2 && pixel_y < 7) || (pixel_x == 216 && pixel_y >= 2 && pixel_y < 8) || (pixel_x == 223 && pixel_y >= 2 && pixel_y < 7) || (pixel_x >= 239 && pixel_x < 241 && pixel_y >= 2 && pixel_y < 4) || (pixel_x == 242 && pixel_y >= 2 && pixel_y < 4) || (pixel_x == 247 && pixel_y >= 2 && pixel_y < 4) || (pixel_x == 250 && pixel_y >= 2 && pixel_y < 7) || (pixel_x == 252 && pixel_y >= 2 && pixel_y < 8) || (pixel_x == 255 && pixel_y >= 2 && pixel_y < 5) || (pixel_x == 258 && pixel_y == 2) || (pixel_x == 261 && pixel_y >= 2 && pixel_y < 7) || (pixel_x == 263 && pixel_y >= 2 && pixel_y < 8) || (pixel_x == 266 && pixel_y >= 2 && pixel_y < 4) || (pixel_x == 268 && pixel_y == 2) || (pixel_x == 275 && pixel_y >= 2 && pixel_y < 8) || (pixel_x == 287 && pixel_y >= 2 && pixel_y < 6) || (pixel_x == 289 && pixel_y >= 2 && pixel_y < 4) || (pixel_x == 293 && pixel_y >= 2 && pixel_y < 7) || (pixel_x == 296 && pixel_y >= 2 && pixel_y < 6) || (pixel_x == 301 && pixel_y >= 2 && pixel_y < 4) || (pixel_x == 303 && pixel_y >= 2 && pixel_y < 4) || (pixel_x >= 308 && pixel_x < 310 && pixel_y == 2) || (pixel_x == 317 && pixel_y >= 2 && pixel_y < 4) || (pixel_x >= 328 && pixel_x < 330 && pixel_y == 2) || (pixel_x == 371 && pixel_y >= 2 && pixel_y < 8) || (pixel_x == 446 && pixel_y >= 2 && pixel_y < 8) || (pixel_x == 484 && pixel_y >= 2 && pixel_y < 9) || (pixel_x == 495 && pixel_y == 2) || (pixel_x == 11 && pixel_y == 3) || (pixel_x == 13 && pixel_y == 3) || (pixel_x == 18 && pixel_y >= 3 && pixel_y < 5) || (pixel_x >= 22 && pixel_x < 25 && pixel_y == 3) || (pixel_x == 28 && pixel_y >= 3 && pixel_y < 5) || (pixel_x == 38 && pixel_y >= 3 && pixel_y < 7) || (pixel_x == 46 && pixel_y >= 3 && pixel_y < 8) || (pixel_x == 83 && pixel_y == 3) || (pixel_x == 88 && pixel_y >= 3 && pixel_y < 8) || (pixel_x == 94 && pixel_y == 3) || (pixel_x == 99 && pixel_y >= 3 && pixel_y < 5) || (pixel_x == 103 && pixel_y == 3) || (pixel_x == 105 && pixel_y >= 3 && pixel_y < 8) || (pixel_x == 109 && pixel_y >= 3 && pixel_y < 5) || (pixel_x == 121 && pixel_y == 3) || (pixel_x >= 125 && pixel_x < 127 && pixel_y >= 3 && pixel_y < 5) || (pixel_x == 136 && pixel_y == 3) || (pixel_x == 141 && pixel_y == 3) || (pixel_x == 148 && pixel_y == 3) || (pixel_x == 156 && pixel_y == 3) || (pixel_x == 163 && pixel_y >= 3 && pixel_y < 5) || (pixel_x == 167 && pixel_y >= 3 && pixel_y < 6) || (pixel_x == 169 && pixel_y >= 3 && pixel_y < 6) || (pixel_x == 212 && pixel_y >= 3 && pixel_y < 5) || (pixel_x >= 226 && pixel_x < 228 && pixel_y >= 3 && pixel_y < 5) || (pixel_x == 257 && pixel_y >= 3 && pixel_y < 7) || (pixel_x == 269 && pixel_y == 3) || (pixel_x == 285 && pixel_y >= 3 && pixel_y < 7) || (pixel_x == 292 && pixel_y >= 3 && pixel_y < 7) || (pixel_x == 297 && pixel_y >= 3 && pixel_y < 6) || (pixel_x == 302 && pixel_y >= 3 && pixel_y < 8) || (pixel_x == 308 && pixel_y == 3) || (pixel_x == 328 && pixel_y == 3) || (pixel_x >= 344 && pixel_x < 347 && pixel_y == 3) || (pixel_x >= 349 && pixel_x < 352 && pixel_y == 3) || (pixel_x >= 355 && pixel_x < 358 && pixel_y == 3) || (pixel_x >= 360 && pixel_x < 362 && pixel_y == 3) || (pixel_x >= 365 && pixel_x < 368 && pixel_y == 3) || (pixel_x == 370 && pixel_y == 3) || (pixel_x >= 372 && pixel_x < 374 && pixel_y == 3) || (pixel_x >= 376 && pixel_x < 379 && pixel_y == 3) || (pixel_x >= 382 && pixel_x < 384 && pixel_y == 3) || (pixel_x >= 386 && pixel_x < 388 && pixel_y == 3) || (pixel_x >= 392 && pixel_x < 395 && pixel_y == 3) || (pixel_x >= 399 && pixel_x < 401 && pixel_y == 3) || (pixel_x >= 407 && pixel_x < 412 && pixel_y == 3) || (pixel_x >= 413 && pixel_x < 417 && pixel_y == 3) || (pixel_x >= 418 && pixel_x < 422 && pixel_y == 3) || (pixel_x >= 423 && pixel_x < 425 && pixel_y >= 3 && pixel_y < 5) || (pixel_x >= 425 && pixel_x < 427 && pixel_y == 3) || (pixel_x >= 430 && pixel_x < 433 && pixel_y == 3) || (pixel_x >= 435 && pixel_x < 438 && pixel_y == 3) || (pixel_x >= 440 && pixel_x < 443 && pixel_y == 3) || (pixel_x == 445 && pixel_y == 3) || (pixel_x == 447 && pixel_y == 3) || (pixel_x == 450 && pixel_y >= 3 && pixel_y < 7) || (pixel_x == 453 && pixel_y >= 3 && pixel_y < 8) || (pixel_x == 455 && pixel_y == 3) || (pixel_x >= 459 && pixel_x < 461 && pixel_y == 3) || (pixel_x == 462 && pixel_y >= 3 && pixel_y < 5) || (pixel_x >= 466 && pixel_x < 468 && pixel_y == 3) || (pixel_x == 469 && pixel_y == 3) || (pixel_x == 471 && pixel_y == 3) || (pixel_x == 475 && pixel_y >= 3 && pixel_y < 5) || (pixel_x >= 477 && pixel_x < 481 && pixel_y == 3) || (pixel_x == 494 && pixel_y == 3) || (pixel_x == 19 && pixel_y >= 4 && pixel_y < 8) || (pixel_x >= 23 && pixel_x < 25 && pixel_y >= 4 && pixel_y < 6) || (pixel_x == 56 && pixel_y >= 4 && pixel_y < 7) || (pixel_x == 77 && pixel_y == 4) || (pixel_x == 80 && pixel_y == 4) || (pixel_x == 93 && pixel_y == 4) || (pixel_x == 98 && pixel_y == 4) || (pixel_x == 102 && pixel_y >= 4 && pixel_y < 6) || (pixel_x == 110 && pixel_y == 4) || (pixel_x == 114 && pixel_y == 4) || (pixel_x == 116 && pixel_y == 4) || (pixel_x == 120 && pixel_y >= 4 && pixel_y < 6) || (pixel_x >= 130 && pixel_x < 132 && pixel_y == 4) || (pixel_x == 147 && pixel_y == 4) || (pixel_x == 151 && pixel_y == 4) || (pixel_x == 153 && pixel_y == 4) || (pixel_x == 157 && pixel_y == 4) || (pixel_x == 172 && pixel_y >= 4 && pixel_y < 7) || (pixel_x == 175 && pixel_y >= 4 && pixel_y < 8) || (pixel_x >= 178 && pixel_x < 180 && pixel_y == 4) || (pixel_x == 182 && pixel_y == 4) || (pixel_x >= 195 && pixel_x < 197 && pixel_y == 4) || (pixel_x >= 200 && pixel_x < 202 && pixel_y == 4) || (pixel_x == 207 && pixel_y >= 4 && pixel_y < 8) || (pixel_x >= 210 && pixel_x < 212 && pixel_y == 4) || (pixel_x == 237 && pixel_y >= 4 && pixel_y < 6) || (pixel_x == 239 && pixel_y == 4) || (pixel_x == 243 && pixel_y == 4) || (pixel_x == 246 && pixel_y == 4) || (pixel_x >= 253 && pixel_x < 255 && pixel_y == 4) || (pixel_x >= 264 && pixel_x < 266 && pixel_y == 4) || (pixel_x == 270 && pixel_y == 4) || (pixel_x == 290 && pixel_y >= 4 && pixel_y < 8) || (pixel_x == 307 && pixel_y >= 4 && pixel_y < 6) || (pixel_x == 318 && pixel_y == 4) || (pixel_x == 327 && pixel_y >= 4 && pixel_y < 6) || (pixel_x == 330 && pixel_y == 4) || (pixel_x == 343 && pixel_y >= 4 && pixel_y < 7) || (pixel_x == 346 && pixel_y >= 4 && pixel_y < 8) || (pixel_x >= 348 && pixel_x < 350 && pixel_y == 4) || (pixel_x == 352 && pixel_y >= 4 && pixel_y < 6) || (pixel_x == 354 && pixel_y >= 4 && pixel_y < 7) || (pixel_x == 359 && pixel_y >= 4 && pixel_y < 7) || (pixel_x == 365 && pixel_y >= 4 && pixel_y < 8) || (pixel_x == 368 && pixel_y == 4) || (pixel_x == 375 && pixel_y >= 4 && pixel_y < 7) || (pixel_x == 378 && pixel_y >= 4 && pixel_y < 10) || (pixel_x == 384 && pixel_y >= 4 && pixel_y < 8) || (pixel_x == 387 && pixel_y >= 4 && pixel_y < 8) || (pixel_x == 394 && pixel_y >= 4 && pixel_y < 9) || (pixel_x >= 398 && pixel_x < 400 && pixel_y == 4) || (pixel_x == 407 && pixel_y >= 4 && pixel_y < 8) || (pixel_x == 409 && pixel_y >= 4 && pixel_y < 8) || (pixel_x == 411 && pixel_y >= 4 && pixel_y < 7) || (pixel_x == 413 && pixel_y >= 4 && pixel_y < 8) || (pixel_x == 416 && pixel_y >= 4 && pixel_y < 8) || (pixel_x == 418 && pixel_y >= 4 && pixel_y < 7) || (pixel_x == 421 && pixel_y >= 4 && pixel_y < 8) || (pixel_x == 427 && pixel_y >= 4 && pixel_y < 6) || (pixel_x == 429 && pixel_y >= 4 && pixel_y < 8) || (pixel_x == 432 && pixel_y >= 4 && pixel_y < 10) || (pixel_x >= 434 && pixel_x < 436 && pixel_y >= 4 && pixel_y < 7) || (pixel_x == 440 && pixel_y == 4) || (pixel_x == 456 && pixel_y >= 4 && pixel_y < 6) || (pixel_x == 463 && pixel_y >= 4 && pixel_y < 6) || (pixel_x >= 467 && pixel_x < 469 && pixel_y >= 4 && pixel_y < 6) || (pixel_x == 472 && pixel_y >= 4 && pixel_y < 6) || (pixel_x == 479 && pixel_y == 4) || (pixel_x == 483 && pixel_y >= 4 && pixel_y < 6) || (pixel_x == 495 && pixel_y >= 4 && pixel_y < 6) || (pixel_x == 11 && pixel_y >= 5 && pixel_y < 7) || (pixel_x == 13 && pixel_y >= 5 && pixel_y < 7) || (pixel_x == 20 && pixel_y >= 5 && pixel_y < 7) || (pixel_x >= 26 && pixel_x < 28 && pixel_y >= 5 && pixel_y < 7) || (pixel_x >= 29 && pixel_x < 31 && pixel_y == 5) || (pixel_x >= 54 && pixel_x < 56 && pixel_y == 5) || (pixel_x == 57 && pixel_y == 5) || (pixel_x >= 81 && pixel_x < 83 && pixel_y == 5) || (pixel_x == 92 && pixel_y >= 5 && pixel_y < 8) || (pixel_x == 100 && pixel_y >= 5 && pixel_y < 7) || (pixel_x >= 103 && pixel_x < 105 && pixel_y == 5) || (pixel_x == 111 && pixel_y >= 5 && pixel_y < 7) || (pixel_x == 119 && pixel_y >= 5 && pixel_y < 8) || (pixel_x == 124 && pixel_y >= 5 && pixel_y < 8) || (pixel_x == 127 && pixel_y >= 5 && pixel_y < 7) || (pixel_x >= 145 && pixel_x < 147 && pixel_y == 5) || (pixel_x >= 158 && pixel_x < 160 && pixel_y == 5) || (pixel_x == 162 && pixel_y == 5) || (pixel_x == 168 && pixel_y == 5) || (pixel_x == 170 && pixel_y == 5) || (pixel_x == 174 && pixel_y == 5) || (pixel_x == 183 && pixel_y >= 5 && pixel_y < 7) || (pixel_x == 227 && pixel_y == 5) || (pixel_x == 238 && pixel_y == 5) || (pixel_x == 240 && pixel_y >= 5 && pixel_y < 7) || (pixel_x == 244 && pixel_y >= 5 && pixel_y < 7) || (pixel_x == 247 && pixel_y >= 5 && pixel_y < 8) || (pixel_x == 253 && pixel_y == 5) || (pixel_x == 265 && pixel_y >= 5 && pixel_y < 7) || (pixel_x == 271 && pixel_y >= 5 && pixel_y < 8) || (pixel_x == 286 && pixel_y >= 5 && pixel_y < 8) || (pixel_x == 306 && pixel_y >= 5 && pixel_y < 8) || (pixel_x == 319 && pixel_y >= 5 && pixel_y < 7) || (pixel_x == 348 && pixel_y >= 5 && pixel_y < 7) || (pixel_x == 367 && pixel_y == 5) || (pixel_x == 398 && pixel_y == 5) || (pixel_x == 423 && pixel_y >= 5 && pixel_y < 10) || (pixel_x >= 441 && pixel_x < 443 && pixel_y == 5) || (pixel_x == 458 && pixel_y >= 5 && pixel_y < 7) || (pixel_x == 461 && pixel_y >= 5 && pixel_y < 8) || (pixel_x == 464 && pixel_y >= 5 && pixel_y < 8) || (pixel_x == 474 && pixel_y >= 5 && pixel_y < 7) || (pixel_x == 478 && pixel_y >= 5 && pixel_y < 8) || (pixel_x == 498 && pixel_y == 5) || (pixel_x >= 500 && pixel_x < 503 && pixel_y == 5) || (pixel_x == 22 && pixel_y >= 6 && pixel_y < 8) || (pixel_x == 24 && pixel_y == 6) || (pixel_x == 30 && pixel_y >= 6 && pixel_y < 8) || (pixel_x == 76 && pixel_y == 6) || (pixel_x == 81 && pixel_y == 6) || (pixel_x == 116 && pixel_y >= 6 && pixel_y < 8) || (pixel_x >= 147 && pixel_x < 149 && pixel_y == 6) || (pixel_x >= 156 && pixel_x < 158 && pixel_y == 6) || (pixel_x == 222 && pixel_y >= 6 && pixel_y < 8) || (pixel_x == 228 && pixel_y == 6) || (pixel_x == 245 && pixel_y >= 6 && pixel_y < 8) || (pixel_x == 258 && pixel_y >= 6 && pixel_y < 8) || (pixel_x == 266 && pixel_y >= 6 && pixel_y < 8) || (pixel_x == 295 && pixel_y >= 6 && pixel_y < 8) || (pixel_x == 298 && pixel_y >= 6 && pixel_y < 8) || (pixel_x == 351 && pixel_y >= 6 && pixel_y < 8) || (pixel_x == 399 && pixel_y == 6) || (pixel_x == 426 && pixel_y >= 6 && pixel_y < 8) || (pixel_x == 431 && pixel_y >= 6 && pixel_y < 8) || (pixel_x >= 442 && pixel_x < 444 && pixel_y == 6) || (pixel_x == 457 && pixel_y >= 6 && pixel_y < 8) || (pixel_x == 467 && pixel_y == 6) || (pixel_x == 469 && pixel_y >= 6 && pixel_y < 8) || (pixel_x == 473 && pixel_y >= 6 && pixel_y < 9) || (pixel_x == 477 && pixel_y >= 6 && pixel_y < 8) || (pixel_x == 494 && pixel_y >= 6 && pixel_y < 9) || (pixel_x == 2 && pixel_y == 7) || (pixel_x >= 17 && pixel_x < 19 && pixel_y == 7) || (pixel_x == 25 && pixel_y == 7) || (pixel_x >= 27 && pixel_x < 30 && pixel_y == 7) || (pixel_x == 31 && pixel_y == 7) || (pixel_x == 39 && pixel_y == 7) || (pixel_x == 61 && pixel_y >= 7 && pixel_y < 9) || (pixel_x == 72 && pixel_y == 7) || (pixel_x == 75 && pixel_y == 7) || (pixel_x >= 82 && pixel_x < 84 && pixel_y == 7) || (pixel_x == 87 && pixel_y == 7) || (pixel_x == 89 && pixel_y == 7) || (pixel_x >= 93 && pixel_x < 95 && pixel_y == 7) || (pixel_x >= 97 && pixel_x < 100 && pixel_y == 7) || (pixel_x >= 108 && pixel_x < 111 && pixel_y == 7) || (pixel_x >= 114 && pixel_x < 116 && pixel_y == 7) || (pixel_x >= 125 && pixel_x < 127 && pixel_y == 7) || (pixel_x >= 129 && pixel_x < 132 && pixel_y == 7) || (pixel_x == 136 && pixel_y == 7) || (pixel_x >= 141 && pixel_x < 143 && pixel_y == 7) || (pixel_x == 156 && pixel_y == 7) || (pixel_x == 162 && pixel_y == 7) || (pixel_x == 167 && pixel_y == 7) || (pixel_x >= 178 && pixel_x < 180 && pixel_y == 7) || (pixel_x >= 184 && pixel_x < 186 && pixel_y == 7) || (pixel_x >= 189 && pixel_x < 191 && pixel_y == 7) || (pixel_x >= 195 && pixel_x < 197 && pixel_y == 7) || (pixel_x >= 205 && pixel_x < 207 && pixel_y == 7) || (pixel_x == 215 && pixel_y == 7) || (pixel_x == 217 && pixel_y == 7) || (pixel_x >= 220 && pixel_x < 222 && pixel_y == 7) || (pixel_x == 229 && pixel_y == 7) || (pixel_x >= 232 && pixel_x < 234 && pixel_y == 7) || (pixel_x >= 248 && pixel_x < 250 && pixel_y == 7) || (pixel_x >= 259 && pixel_x < 261 && pixel_y == 7) || (pixel_x >= 269 && pixel_x < 271 && pixel_y == 7) || (pixel_x >= 280 && pixel_x < 282 && pixel_y == 7) || (pixel_x >= 307 && pixel_x < 310 && pixel_y == 7) || (pixel_x == 320 && pixel_y == 7) || (pixel_x >= 344 && pixel_x < 346 && pixel_y == 7) || (pixel_x >= 349 && pixel_x < 351 && pixel_y == 7) || (pixel_x >= 355 && pixel_x < 358 && pixel_y == 7) || (pixel_x >= 360 && pixel_x < 362 && pixel_y == 7) || (pixel_x >= 366 && pixel_x < 368 && pixel_y == 7) || (pixel_x >= 376 && pixel_x < 378 && pixel_y == 7) || (pixel_x == 388 && pixel_y == 7) || (pixel_x == 400 && pixel_y == 7) || (pixel_x == 404 && pixel_y == 7) || (pixel_x >= 419 && pixel_x < 421 && pixel_y == 7) || (pixel_x >= 424 && pixel_x < 426 && pixel_y == 7) || (pixel_x == 430 && pixel_y == 7) || (pixel_x >= 440 && pixel_x < 443 && pixel_y == 7) || (pixel_x >= 447 && pixel_x < 449 && pixel_y == 7) || (pixel_x >= 451 && pixel_x < 453 && pixel_y == 7) || (pixel_x == 466 && pixel_y == 7) || (pixel_x >= 479 && pixel_x < 481 && pixel_y == 7) || (pixel_x == 40 && pixel_y == 8) || (pixel_x >= 44 && pixel_x < 46 && pixel_y == 8) || (pixel_x == 142 && pixel_y == 8) || (pixel_x == 260 && pixel_y == 8) || (pixel_x >= 332 && pixel_x < 336 && pixel_y == 8) || (pixel_x == 141 && pixel_y == 9) || (pixel_x == 261 && pixel_y == 9) || (pixel_x >= 313 && pixel_x < 315 && pixel_y == 9) || (pixel_x >= 322 && pixel_x < 324 && pixel_y == 9) || (pixel_x >= 375 && pixel_x < 378 && pixel_y == 9) || (pixel_x >= 392 && pixel_x < 394 && pixel_y == 9) || (pixel_x >= 471 && pixel_x < 473 && pixel_y == 9) || (pixel_x == 485 && pixel_y == 9) || (pixel_x == 493 && pixel_y == 9))
    hit <= 1;
else hit <= 0;

endmodule
