module registerRenderer (
  input [10:0] x, y,
  input [2:0] r, g, b,
  input [3:0] registerIndex,
  input [15:0] registerValue
);

endmodule
